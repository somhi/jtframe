/*  This file is part of JTFRAME.
    JTFRAME program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JTFRAME program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JTFRAME.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 7-3-2019 */

module jtframe_led(
    input        rst,
    input        clk,
    input        LVBL,
    input        downloading,
    input        osd_shown,
    input [3:0]  gfx_en,
    input [7:0]  debug_bus,
    input [1:0]  game_led,
    input        cheat_led,
    output reg   led
);

wire  sys_led, enlarged, debug_led;
reg   last_LVBL, cen_VB;

`ifdef MISTER
localparam POL = 1;
`else
localparam POL = 0;
`endif

`ifdef JTFRAME_DEBUG
    reg [6:0] fcnt;
    always @(posedge clk,posedge rst) begin
        if( rst ) begin
            fcnt <= 0;
        end else begin
            if( !LVBL && last_LVBL ) fcnt <= fcnt+1;
        end
    end
    assign debug_led = debug_bus==0 && fcnt[6];
`else
    assign debug_led = 0;
`endif

// debug_led is XOR'ed because it blinks
assign sys_led = ~( downloading | cheat_led /*| osd_shown*/ | (|(~gfx_en)))^debug_led;

always @(posedge clk) begin
    last_LVBL <= LVBL;
    cen_VB    <= !LVBL && last_LVBL;
end

// Make the minimum pulse length equal to 16 frames = 0.26s
jtframe_enlarger #(.W(4)) u_enlarger(
    .rst        ( rst               ),
    .clk        ( clk               ),
    .cen        ( cen_VB            ),
    .pulse_in   ( game_led[0]       ),
    .pulse_out  ( enlarged          )
);

///////////////// LED is on while
// downloading, PLL lock lost, OSD is shown or in reset state
always @(posedge clk, posedge rst) begin
    if( rst ) begin
        led <= POL[0];
    end else begin
        led <= (~enlarged & sys_led ) ^ POL[0];
    end
end

endmodule