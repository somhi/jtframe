// Translation to verilog of Oregano's 8051 core

module addsub_ovcy_4
  (input  [3:0] opa_i,
   input  [3:0] opb_i,
   input  addsub_i,
   input  cy_i,
   output cy_o,
   output ov_o,
   output [3:0] rslt_o);
  wire [2:0] n11190_o;
  wire [2:0] n11191_o;
  wire n11192_o;
  wire n11193_o;
  wire [3:0] n11195_o;
  wire [4:0] n11196_o;
  wire [3:0] n11197_o;
  wire [4:0] n11198_o;
  wire [4:0] n11199_o;
  wire n11201_o;
  wire [1:0] n11202_o;
  wire [2:0] n11203_o;
  wire [1:0] n11204_o;
  wire [2:0] n11205_o;
  wire [2:0] n11206_o;
  wire [3:0] n11208_o;
  wire [4:0] n11209_o;
  wire [3:0] n11210_o;
  wire [4:0] n11211_o;
  wire [4:0] n11212_o;
  wire n11214_o;
  wire [1:0] n11215_o;
  wire [2:0] n11216_o;
  wire [1:0] n11217_o;
  wire [2:0] n11218_o;
  wire [2:0] n11219_o;
  wire [4:0] n11221_o;
  wire [2:0] n11224_o;
  wire n11225_o;
  wire n11226_o;
  wire n11227_o;
  wire n11228_o;
  wire n11229_o;
  wire n11230_o;
  wire n11231_o;
  wire n11232_o;
  wire n11233_o;
  wire n11234_o;
  wire [2:0] n11235_o;
  wire n11236_o;
  wire [3:0] n11242_o;
  assign cy_o = n11225_o;
  assign ov_o = n11234_o;
  assign rslt_o = n11242_o;
  /* addsub_ovcy_rtl.vhd:111:47  */
  assign n11190_o = opa_i[2:0];
  /* addsub_ovcy_rtl.vhd:112:47  */
  assign n11191_o = opb_i[2:0];
  /* addsub_ovcy_rtl.vhd:113:23  */
  assign n11192_o = opa_i[3];
  /* addsub_ovcy_rtl.vhd:114:23  */
  assign n11193_o = opb_i[3];
  assign n11195_o = {n11190_o, 1'b1};
  /* addsub_ovcy_rtl.vhd:118:21  */
  assign n11196_o = {1'b0, n11195_o};  //  uext
  assign n11197_o = {n11191_o, cy_i};
  /* addsub_ovcy_rtl.vhd:118:49  */
  assign n11198_o = {1'b0, n11197_o};  //  uext
  /* addsub_ovcy_rtl.vhd:118:49  */
  assign n11199_o = n11196_o + n11198_o;
  /* addsub_ovcy_rtl.vhd:120:28  */
  assign n11201_o = n11199_o[4];
  assign n11202_o = {n11192_o, 1'b1};
  /* addsub_ovcy_rtl.vhd:121:22  */
  assign n11203_o = {1'b0, n11202_o};  //  uext
  assign n11204_o = {n11193_o, n11201_o};
  /* addsub_ovcy_rtl.vhd:121:44  */
  assign n11205_o = {1'b0, n11204_o};  //  uext
  /* addsub_ovcy_rtl.vhd:121:44  */
  assign n11206_o = n11203_o + n11205_o;
  assign n11208_o = {n11190_o, 1'b0};
  /* addsub_ovcy_rtl.vhd:125:21  */
  assign n11209_o = {1'b0, n11208_o};  //  uext
  assign n11210_o = {n11191_o, cy_i};
  /* addsub_ovcy_rtl.vhd:125:49  */
  assign n11211_o = {1'b0, n11210_o};  //  uext
  /* addsub_ovcy_rtl.vhd:125:49  */
  assign n11212_o = n11209_o - n11211_o;
  /* addsub_ovcy_rtl.vhd:127:28  */
  assign n11214_o = n11212_o[4];
  assign n11215_o = {n11192_o, 1'b0};
  /* addsub_ovcy_rtl.vhd:128:22  */
  assign n11216_o = {1'b0, n11215_o};  //  uext
  assign n11217_o = {n11193_o, n11214_o};
  /* addsub_ovcy_rtl.vhd:128:44  */
  assign n11218_o = {1'b0, n11217_o};  //  uext
  /* addsub_ovcy_rtl.vhd:128:44  */
  assign n11219_o = n11216_o - n11218_o;
  /* addsub_ovcy_rtl.vhd:115:7  */
  assign n11221_o = addsub_i ? n11199_o : n11212_o;
  /* addsub_ovcy_rtl.vhd:115:7  */
  assign n11224_o = addsub_i ? n11206_o : n11219_o;
  /* addsub_ovcy_rtl.vhd:130:24  */
  assign n11225_o = n11224_o[2];
  /* addsub_ovcy_rtl.vhd:131:24  */
  assign n11226_o = n11221_o[4];
  /* addsub_ovcy_rtl.vhd:131:50  */
  assign n11227_o = n11224_o[2];
  /* addsub_ovcy_rtl.vhd:131:37  */
  assign n11228_o = ~n11227_o;
  /* addsub_ovcy_rtl.vhd:131:33  */
  assign n11229_o = n11226_o & n11228_o;
  /* addsub_ovcy_rtl.vhd:132:23  */
  assign n11230_o = n11224_o[2];
  /* addsub_ovcy_rtl.vhd:132:43  */
  assign n11231_o = n11221_o[4];
  /* addsub_ovcy_rtl.vhd:132:31  */
  assign n11232_o = ~n11231_o;
  /* addsub_ovcy_rtl.vhd:132:27  */
  assign n11233_o = n11230_o & n11232_o;
  /* addsub_ovcy_rtl.vhd:131:56  */
  assign n11234_o = n11229_o | n11233_o;
  /* addsub_ovcy_rtl.vhd:133:44  */
  assign n11235_o = n11221_o[3:1];
  /* addsub_ovcy_rtl.vhd:134:36  */
  assign n11236_o = n11224_o[1];
  assign n11242_o = {n11236_o, n11235_o};
endmodule

module addsub_cy_4
  (input  [3:0] opa_i,
   input  [3:0] opb_i,
   input  addsub_i,
   input  cy_i,
   output cy_o,
   output [3:0] rslt_o);
  wire [4:0] n11162_o;
  wire [5:0] n11163_o;
  wire [4:0] n11164_o;
  wire [5:0] n11165_o;
  wire [5:0] n11166_o;
  wire [4:0] n11168_o;
  wire [5:0] n11169_o;
  wire [4:0] n11170_o;
  wire [5:0] n11171_o;
  wire [5:0] n11172_o;
  wire [5:0] n11174_o;
  wire n11175_o;
  wire [3:0] n11176_o;
  assign cy_o = n11175_o;
  assign rslt_o = n11176_o;
  assign n11162_o = {opa_i, 1'b1};
  /* addsub_cy_rtl.vhd:84:19  */
  assign n11163_o = {1'b0, n11162_o};  //  uext
  /* dcml_adjust_rtl.vhd:76:14  */
  assign n11164_o = {opb_i, cy_i};
  /* addsub_cy_rtl.vhd:84:47  */
  assign n11165_o = {1'b0, n11164_o};  //  uext
  /* addsub_cy_rtl.vhd:84:47  */
  assign n11166_o = n11163_o + n11165_o;
  /* dcml_adjust_rtl.vhd:74:14  */
  assign n11168_o = {opa_i, 1'b0};
  /* addsub_cy_rtl.vhd:88:19  */
  assign n11169_o = {1'b0, n11168_o};  //  uext
  /* dcml_adjust_rtl.vhd:73:14  */
  assign n11170_o = {opb_i, cy_i};
  /* addsub_cy_rtl.vhd:88:47  */
  assign n11171_o = {1'b0, n11170_o};  //  uext
  /* addsub_cy_rtl.vhd:88:47  */
  assign n11172_o = n11169_o - n11171_o;
  /* addsub_cy_rtl.vhd:81:5  */
  assign n11174_o = addsub_i ? n11166_o : n11172_o;
  /* addsub_cy_rtl.vhd:90:21  */
  assign n11175_o = n11174_o[5];
  /* addsub_cy_rtl.vhd:91:23  */
  assign n11176_o = n11174_o[4:1];
endmodule

module dcml_adjust_8
  (input  [7:0] data_i,
   input  [1:0] cy_i,
   output [7:0] data_o,
   output cy_o);
  wire [8:0] n11085_o;
  wire [3:0] n11086_o;
  wire n11087_o;
  wire n11089_o;
  wire n11090_o;
  wire [8:0] n11091_o;
  wire [3:0] n11092_o;
  wire [4:0] n11093_o;
  wire [4:0] n11095_o;
  wire n11096_o;
  wire [3:0] n11097_o;
  wire n11098_o;
  wire n11099_o;
  wire n11100_o;
  wire [3:0] n11101_o;
  wire [8:0] n11102_o;
  wire [3:0] n11103_o;
  wire [4:0] n11104_o;
  wire [4:0] n11105_o;
  wire [4:0] n11106_o;
  wire [8:0] n11107_o;
  wire n11108_o;
  wire n11109_o;
  wire [1:0] n11110_o;
  wire n11111_o;
  wire n11112_o;
  wire [1:0] n11113_o;
  wire [1:0] n11114_o;
  wire [8:0] n11118_o;
  wire [8:0] n11119_o;
  wire [8:0] n11120_o;
  wire [3:0] n11124_o;
  wire n11126_o;
  wire n11128_o;
  wire n11129_o;
  wire [3:0] n11130_o;
  wire [4:0] n11131_o;
  wire [4:0] n11133_o;
  wire [4:0] n11134_o;
  wire [4:0] n11135_o;
  wire [4:0] n11136_o;
  wire [4:0] n11137_o;
  wire [3:0] n11138_o;
  wire [3:0] n11139_o;
  wire [3:0] n11140_o;
  wire [8:0] n11141_o;
  wire n11142_o;
  wire n11143_o;
  wire n11144_o;
  wire n11145_o;
  wire n11146_o;
  wire n11147_o;
  wire [1:0] n11148_o;
  wire n11149_o;
  wire [8:0] n11150_o;
  wire [7:0] n11151_o;
  assign data_o = n11151_o;
  assign cy_o = n11149_o;
  /* comb_divider_rtl.vhd:103:47  */
  assign n11085_o = {1'b0, data_i};
  /* dcml_adjust_rtl.vhd:101:28  */
  assign n11086_o = n11085_o[3:0];
  /* dcml_adjust_rtl.vhd:103:17  */
  assign n11087_o = cy_i[0];
  /* dcml_adjust_rtl.vhd:103:41  */
  assign n11089_o = $unsigned(n11086_o) > $unsigned(4'b1001);
  /* dcml_adjust_rtl.vhd:103:28  */
  assign n11090_o = n11087_o | n11089_o;
  /* comb_divider_rtl.vhd:88:7  */
  assign n11091_o = {1'b0, data_i};
  /* dcml_adjust_rtl.vhd:109:36  */
  assign n11092_o = n11091_o[3:0];
  /* dcml_adjust_rtl.vhd:109:55  */
  assign n11093_o = {1'b0, n11092_o};  //  uext
  /* dcml_adjust_rtl.vhd:109:55  */
  assign n11095_o = n11093_o + 5'b00110;
  /* dcml_adjust_rtl.vhd:111:36  */
  assign n11096_o = n11095_o[4];
  /* dcml_adjust_rtl.vhd:112:54  */
  assign n11097_o = n11095_o[3:0];
  /* dcml_adjust_rtl.vhd:120:34  */
  assign n11098_o = n11095_o[4];
  /* dcml_adjust_rtl.vhd:120:45  */
  assign n11099_o = cy_i[0];
  /* dcml_adjust_rtl.vhd:120:38  */
  assign n11100_o = n11098_o | n11099_o;
  /* comb_divider_rtl.vhd:103:47  */
  assign n11101_o = data_i[7:4];
  /* comb_divider_rtl.vhd:75:3  */
  assign n11102_o = {1'b0, n11101_o, n11097_o};
  /* dcml_adjust_rtl.vhd:127:54  */
  assign n11103_o = n11102_o[7:4];
  /* dcml_adjust_rtl.vhd:128:22  */
  assign n11104_o = {4'b0, n11096_o};  //  uext
  /* dcml_adjust_rtl.vhd:127:76  */
  assign n11105_o = {1'b0, n11103_o};  //  uext
  /* dcml_adjust_rtl.vhd:127:76  */
  assign n11106_o = n11105_o + n11104_o;
  /* comb_divider_rtl.vhd:77:14  */
  assign n11107_o = {n11106_o, n11097_o};
  /* dcml_adjust_rtl.vhd:131:33  */
  assign n11108_o = n11107_o[8];
  assign n11109_o = cy_i[1];
  assign n11110_o = {n11109_o, n11100_o};
  /* dcml_adjust_rtl.vhd:131:49  */
  assign n11111_o = n11110_o[1];
  /* dcml_adjust_rtl.vhd:131:42  */
  assign n11112_o = n11108_o | n11111_o;
  assign n11113_o = {n11112_o, n11100_o};
  /* dcml_adjust_rtl.vhd:103:9  */
  assign n11114_o = n11090_o ? n11113_o : cy_i;
  assign n11118_o = {n11106_o, n11097_o};
  assign n11119_o = {1'b0, data_i};
  /* dcml_adjust_rtl.vhd:103:9  */
  assign n11120_o = n11090_o ? n11118_o : n11119_o;
  /* dcml_adjust_rtl.vhd:87:51  */
  assign n11124_o = n11120_o[7:4];
  /* dcml_adjust_rtl.vhd:88:17  */
  assign n11126_o = n11114_o[1];
  /* dcml_adjust_rtl.vhd:88:41  */
  assign n11128_o = $unsigned(n11124_o) > $unsigned(4'b1001);
  /* dcml_adjust_rtl.vhd:88:28  */
  assign n11129_o = n11126_o | n11128_o;
  /* dcml_adjust_rtl.vhd:90:50  */
  assign n11130_o = n11120_o[7:4];
  /* dcml_adjust_rtl.vhd:90:72  */
  assign n11131_o = {1'b0, n11130_o};  //  uext
  /* dcml_adjust_rtl.vhd:90:72  */
  assign n11133_o = n11131_o + 5'b00110;
  assign n11134_o = n11118_o[8:4];
  assign n11135_o = n11119_o[8:4];
  /* dcml_adjust_rtl.vhd:103:9  */
  assign n11136_o = n11090_o ? n11134_o : n11135_o;
  /* dcml_adjust_rtl.vhd:88:9  */
  assign n11137_o = n11129_o ? n11133_o : n11136_o;
  assign n11138_o = n11118_o[3:0];
  assign n11139_o = n11119_o[3:0];
  /* dcml_adjust_rtl.vhd:103:9  */
  assign n11140_o = n11090_o ? n11138_o : n11139_o;
  assign n11141_o = {n11137_o, n11140_o};
  /* dcml_adjust_rtl.vhd:98:27  */
  assign n11142_o = n11141_o[8];
  /* dcml_adjust_rtl.vhd:98:43  */
  assign n11143_o = n11114_o[1];
  /* dcml_adjust_rtl.vhd:98:36  */
  assign n11144_o = n11142_o | n11143_o;
  assign n11145_o = n11113_o[0];
  assign n11146_o = cy_i[0];
  /* dcml_adjust_rtl.vhd:103:9  */
  assign n11147_o = n11090_o ? n11145_o : n11146_o;
  assign n11148_o = {n11144_o, n11147_o};
  /* dcml_adjust_rtl.vhd:138:17  */
  assign n11149_o = n11148_o[1];
  assign n11150_o = {n11137_o, n11140_o};
  /* dcml_adjust_rtl.vhd:139:39  */
  assign n11151_o = n11150_o[7:0];
endmodule

module comb_divider_8
  (input  [7:0] dvdnd_i,
   input  [7:0] dvsor_i,
   output [7:0] qutnt_o,
   output [7:0] rmndr_o);
  wire n10918_o;
  wire [7:0] n10919_o;
  wire n10920_o;
  wire n10922_o;
  wire [7:0] n10923_o;
  wire [7:0] n10924_o;
  wire n10925_o;
  wire n10926_o;
  wire [1:0] n10930_o;
  wire [1:0] n10931_o;
  wire [1:0] n10932_o;
  wire [5:0] n10933_o;
  wire n10935_o;
  wire [7:0] n10936_o;
  wire [1:0] n10937_o;
  wire [7:0] n10938_o;
  wire n10939_o;
  wire [7:0] n10941_o;
  wire [1:0] n10942_o;
  wire [7:0] n10943_o;
  wire [7:0] n10944_o;
  wire [1:0] n10945_o;
  wire n10946_o;
  wire [2:0] n10951_o;
  wire n10952_o;
  wire [2:0] n10953_o;
  wire [2:0] n10954_o;
  wire [4:0] n10955_o;
  wire n10957_o;
  wire [7:0] n10958_o;
  wire [2:0] n10959_o;
  wire [7:0] n10960_o;
  wire n10961_o;
  wire [7:0] n10963_o;
  wire [2:0] n10964_o;
  wire [7:0] n10965_o;
  wire [7:0] n10966_o;
  wire [2:0] n10967_o;
  wire n10968_o;
  wire [3:0] n10973_o;
  wire n10974_o;
  wire [3:0] n10975_o;
  wire [3:0] n10976_o;
  wire [3:0] n10977_o;
  wire n10979_o;
  wire [7:0] n10980_o;
  wire [3:0] n10981_o;
  wire [7:0] n10982_o;
  wire n10983_o;
  wire [7:0] n10985_o;
  wire [3:0] n10986_o;
  wire [7:0] n10987_o;
  wire [7:0] n10988_o;
  wire [3:0] n10989_o;
  wire n10990_o;
  wire [4:0] n10995_o;
  wire n10996_o;
  wire [4:0] n10997_o;
  wire [4:0] n10998_o;
  wire [2:0] n10999_o;
  wire n11001_o;
  wire [7:0] n11002_o;
  wire [4:0] n11003_o;
  wire [7:0] n11004_o;
  wire n11005_o;
  wire [7:0] n11007_o;
  wire [4:0] n11008_o;
  wire [7:0] n11009_o;
  wire [7:0] n11010_o;
  wire [4:0] n11011_o;
  wire n11012_o;
  wire [5:0] n11017_o;
  wire n11018_o;
  wire [5:0] n11019_o;
  wire [5:0] n11020_o;
  wire [1:0] n11021_o;
  wire n11023_o;
  wire [7:0] n11024_o;
  wire [5:0] n11025_o;
  wire [7:0] n11026_o;
  wire n11027_o;
  wire [7:0] n11029_o;
  wire [5:0] n11030_o;
  wire [7:0] n11031_o;
  wire [7:0] n11032_o;
  wire [5:0] n11033_o;
  wire n11034_o;
  wire [6:0] n11039_o;
  wire n11040_o;
  wire [6:0] n11041_o;
  wire [6:0] n11042_o;
  wire n11043_o;
  wire n11045_o;
  wire [7:0] n11046_o;
  wire [6:0] n11047_o;
  wire [7:0] n11048_o;
  wire n11049_o;
  wire [7:0] n11051_o;
  wire [6:0] n11052_o;
  wire [7:0] n11053_o;
  wire [7:0] n11054_o;
  wire [6:0] n11055_o;
  wire n11056_o;
  wire [7:0] n11061_o;
  wire [7:0] n11062_o;
  wire [7:0] n11063_o;
  wire n11065_o;
  wire n11066_o;
  wire [7:0] n11068_o;
  wire [7:0] n11070_o;
  wire n11071_o;
  wire [7:0] n11072_o;
  assign qutnt_o = n11072_o;
  assign rmndr_o = n11070_o;
  /* comb_divider_rtl.vhd:88:44  */
  assign n10918_o = dvdnd_i[7];
  /* comb_divider_rtl.vhd:88:10  */
  assign n10919_o = {7'b0, n10918_o};  //  uext
  /* comb_divider_rtl.vhd:88:72  */
  assign n10920_o = $unsigned(n10919_o) >= $unsigned(dvsor_i);
  /* comb_divider_rtl.vhd:92:47  */
  assign n10922_o = dvdnd_i[7];
  /* comb_divider_rtl.vhd:92:21  */
  assign n10923_o = {7'b0, n10922_o};  //  uext
  /* comb_divider_rtl.vhd:93:21  */
  assign n10924_o = n10923_o - dvsor_i;
  /* comb_divider_rtl.vhd:97:54  */
  assign n10925_o = n10924_o[0];
  /* comb_divider_rtl.vhd:98:39  */
  assign n10926_o = dvdnd_i[6];
  assign n10930_o = {n10925_o, n10926_o};
  assign n10931_o = dvdnd_i[7:6];
  /* comb_divider_rtl.vhd:88:7  */
  assign n10932_o = n10920_o ? n10930_o : n10931_o;
  assign n10933_o = dvdnd_i[5:0];
  /* comb_divider_rtl.vhd:88:7  */
  assign n10935_o = n10920_o ? 1'b1 : 1'b0;
  assign n10936_o = {n10932_o, n10933_o};
  /* comb_divider_rtl.vhd:88:44  */
  assign n10937_o = n10936_o[7:6];
  /* comb_divider_rtl.vhd:88:10  */
  assign n10938_o = {6'b0, n10937_o};  //  uext
  /* comb_divider_rtl.vhd:88:72  */
  assign n10939_o = $unsigned(n10938_o) >= $unsigned(dvsor_i);
  assign n10941_o = {n10932_o, n10933_o};
  /* comb_divider_rtl.vhd:92:47  */
  assign n10942_o = n10941_o[7:6];
  /* comb_divider_rtl.vhd:92:21  */
  assign n10943_o = {6'b0, n10942_o};  //  uext
  /* comb_divider_rtl.vhd:93:21  */
  assign n10944_o = n10943_o - dvsor_i;
  /* comb_divider_rtl.vhd:97:54  */
  assign n10945_o = n10944_o[1:0];
  /* comb_divider_rtl.vhd:98:39  */
  assign n10946_o = dvdnd_i[5];
  assign n10951_o = {n10945_o, n10946_o};
  assign n10952_o = dvdnd_i[5];
  assign n10953_o = {n10932_o, n10952_o};
  /* comb_divider_rtl.vhd:88:7  */
  assign n10954_o = n10939_o ? n10951_o : n10953_o;
  assign n10955_o = dvdnd_i[4:0];
  /* comb_divider_rtl.vhd:88:7  */
  assign n10957_o = n10939_o ? 1'b1 : 1'b0;
  assign n10958_o = {n10954_o, n10955_o};
  /* comb_divider_rtl.vhd:88:44  */
  assign n10959_o = n10958_o[7:5];
  /* comb_divider_rtl.vhd:88:10  */
  assign n10960_o = {5'b0, n10959_o};  //  uext
  /* comb_divider_rtl.vhd:88:72  */
  assign n10961_o = $unsigned(n10960_o) >= $unsigned(dvsor_i);
  assign n10963_o = {n10954_o, n10955_o};
  /* comb_divider_rtl.vhd:92:47  */
  assign n10964_o = n10963_o[7:5];
  /* comb_divider_rtl.vhd:92:21  */
  assign n10965_o = {5'b0, n10964_o};  //  uext
  /* comb_divider_rtl.vhd:93:21  */
  assign n10966_o = n10965_o - dvsor_i;
  /* comb_divider_rtl.vhd:97:54  */
  assign n10967_o = n10966_o[2:0];
  /* comb_divider_rtl.vhd:98:39  */
  assign n10968_o = dvdnd_i[4];
  assign n10973_o = {n10967_o, n10968_o};
  assign n10974_o = dvdnd_i[4];
  assign n10975_o = {n10954_o, n10974_o};
  /* comb_divider_rtl.vhd:88:7  */
  assign n10976_o = n10961_o ? n10973_o : n10975_o;
  assign n10977_o = dvdnd_i[3:0];
  /* comb_divider_rtl.vhd:88:7  */
  assign n10979_o = n10961_o ? 1'b1 : 1'b0;
  assign n10980_o = {n10976_o, n10977_o};
  /* comb_divider_rtl.vhd:88:44  */
  assign n10981_o = n10980_o[7:4];
  /* comb_divider_rtl.vhd:88:10  */
  assign n10982_o = {4'b0, n10981_o};  //  uext
  /* comb_divider_rtl.vhd:88:72  */
  assign n10983_o = $unsigned(n10982_o) >= $unsigned(dvsor_i);
  assign n10985_o = {n10976_o, n10977_o};
  /* comb_divider_rtl.vhd:92:47  */
  assign n10986_o = n10985_o[7:4];
  /* comb_divider_rtl.vhd:92:21  */
  assign n10987_o = {4'b0, n10986_o};  //  uext
  /* comb_divider_rtl.vhd:93:21  */
  assign n10988_o = n10987_o - dvsor_i;
  /* comb_divider_rtl.vhd:97:54  */
  assign n10989_o = n10988_o[3:0];
  /* comb_divider_rtl.vhd:98:39  */
  assign n10990_o = dvdnd_i[3];
  assign n10995_o = {n10989_o, n10990_o};
  assign n10996_o = dvdnd_i[3];
  assign n10997_o = {n10976_o, n10996_o};
  /* comb_divider_rtl.vhd:88:7  */
  assign n10998_o = n10983_o ? n10995_o : n10997_o;
  assign n10999_o = dvdnd_i[2:0];
  /* comb_divider_rtl.vhd:88:7  */
  assign n11001_o = n10983_o ? 1'b1 : 1'b0;
  assign n11002_o = {n10998_o, n10999_o};
  /* comb_divider_rtl.vhd:88:44  */
  assign n11003_o = n11002_o[7:3];
  /* comb_divider_rtl.vhd:88:10  */
  assign n11004_o = {3'b0, n11003_o};  //  uext
  /* comb_divider_rtl.vhd:88:72  */
  assign n11005_o = $unsigned(n11004_o) >= $unsigned(dvsor_i);
  assign n11007_o = {n10998_o, n10999_o};
  /* comb_divider_rtl.vhd:92:47  */
  assign n11008_o = n11007_o[7:3];
  /* comb_divider_rtl.vhd:92:21  */
  assign n11009_o = {3'b0, n11008_o};  //  uext
  /* comb_divider_rtl.vhd:93:21  */
  assign n11010_o = n11009_o - dvsor_i;
  /* comb_divider_rtl.vhd:97:54  */
  assign n11011_o = n11010_o[4:0];
  /* comb_divider_rtl.vhd:98:39  */
  assign n11012_o = dvdnd_i[2];
  assign n11017_o = {n11011_o, n11012_o};
  assign n11018_o = dvdnd_i[2];
  assign n11019_o = {n10998_o, n11018_o};
  /* comb_divider_rtl.vhd:88:7  */
  assign n11020_o = n11005_o ? n11017_o : n11019_o;
  assign n11021_o = dvdnd_i[1:0];
  /* comb_divider_rtl.vhd:88:7  */
  assign n11023_o = n11005_o ? 1'b1 : 1'b0;
  assign n11024_o = {n11020_o, n11021_o};
  /* comb_divider_rtl.vhd:88:44  */
  assign n11025_o = n11024_o[7:2];
  /* comb_divider_rtl.vhd:88:10  */
  assign n11026_o = {2'b0, n11025_o};  //  uext
  /* comb_divider_rtl.vhd:88:72  */
  assign n11027_o = $unsigned(n11026_o) >= $unsigned(dvsor_i);
  assign n11029_o = {n11020_o, n11021_o};
  /* comb_divider_rtl.vhd:92:47  */
  assign n11030_o = n11029_o[7:2];
  /* comb_divider_rtl.vhd:92:21  */
  assign n11031_o = {2'b0, n11030_o};  //  uext
  /* comb_divider_rtl.vhd:93:21  */
  assign n11032_o = n11031_o - dvsor_i;
  /* comb_divider_rtl.vhd:97:54  */
  assign n11033_o = n11032_o[5:0];
  /* comb_divider_rtl.vhd:98:39  */
  assign n11034_o = dvdnd_i[1];
  assign n11039_o = {n11033_o, n11034_o};
  assign n11040_o = dvdnd_i[1];
  assign n11041_o = {n11020_o, n11040_o};
  /* comb_divider_rtl.vhd:88:7  */
  assign n11042_o = n11027_o ? n11039_o : n11041_o;
  assign n11043_o = dvdnd_i[0];
  /* comb_divider_rtl.vhd:88:7  */
  assign n11045_o = n11027_o ? 1'b1 : 1'b0;
  assign n11046_o = {n11042_o, n11043_o};
  /* comb_divider_rtl.vhd:88:44  */
  assign n11047_o = n11046_o[7:1];
  /* comb_divider_rtl.vhd:88:10  */
  assign n11048_o = {1'b0, n11047_o};  //  uext
  /* comb_divider_rtl.vhd:88:72  */
  assign n11049_o = $unsigned(n11048_o) >= $unsigned(dvsor_i);
  assign n11051_o = {n11042_o, n11043_o};
  /* comb_divider_rtl.vhd:92:47  */
  assign n11052_o = n11051_o[7:1];
  /* comb_divider_rtl.vhd:92:21  */
  assign n11053_o = {1'b0, n11052_o};  //  uext
  /* comb_divider_rtl.vhd:93:21  */
  assign n11054_o = n11053_o - dvsor_i;
  /* comb_divider_rtl.vhd:97:54  */
  assign n11055_o = n11054_o[6:0];
  /* comb_divider_rtl.vhd:98:39  */
  assign n11056_o = dvdnd_i[0];
  assign n11061_o = {n11055_o, n11056_o};
  assign n11062_o = {n11042_o, n11043_o};
  /* comb_divider_rtl.vhd:103:47  */
  assign n11063_o = n11049_o ? n11061_o : n11062_o;
  /* comb_divider_rtl.vhd:88:7  */
  assign n11065_o = n11049_o ? 1'b1 : 1'b0;
  /* comb_divider_rtl.vhd:88:72  */
  assign n11066_o = $unsigned(n11063_o) >= $unsigned(dvsor_i);
  /* comb_divider_rtl.vhd:93:21  */
  assign n11068_o = n11063_o - dvsor_i;
  /* comb_divider_rtl.vhd:88:7  */
  assign n11070_o = n11066_o ? n11068_o : n11063_o;
  /* comb_divider_rtl.vhd:88:7  */
  assign n11071_o = n11066_o ? 1'b1 : 1'b0;
  assign n11072_o = {n10935_o, n10957_o, n10979_o, n11001_o, n11023_o, n11045_o, n11065_o, n11071_o};
endmodule

module comb_mltplr_8
  (input  [7:0] mltplcnd_i,
   input  [7:0] mltplctr_i,
   output [15:0] product_o);
  wire [15:0] n10908_o;
  wire [15:0] n10909_o;
  wire [15:0] n10910_o;
  assign product_o = n10910_o;
  /* comb_mltplr_rtl.vhd:81:32  */
  assign n10908_o = {8'b0, mltplctr_i};  //  uext
  /* comb_mltplr_rtl.vhd:81:32  */
  assign n10909_o = {8'b0, mltplcnd_i};  //  uext
  /* comb_mltplr_rtl.vhd:81:32  */
  assign n10910_o = n10908_o * n10909_o; // umul
endmodule

module addsub_core_8
  (input  [7:0] opa_i,
   input  [7:0] opb_i,
   input  addsub_i,
   input  cy_i,
   output [1:0] cy_o,
   output ov_o,
   output [7:0] rslt_o);
  wire [2:0] s_cy;
  wire [3:0] n10879_o;
  wire [3:0] n10880_o;
  wire n10881_o;
  wire gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_n10882;
  wire [3:0] gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_n10883;
  wire gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_cy_o;
  wire [3:0] gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_rslt_o;
  wire n10888_o;
  wire [3:0] n10889_o;
  wire [3:0] n10890_o;
  wire n10891_o;
  wire gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_n10892;
  wire gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_n10893;
  wire [3:0] gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_n10894;
  wire gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_cy_o;
  wire gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_ov_o;
  wire [3:0] gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_rslt_o;
  wire [2:0] n10902_o;
  wire [1:0] n10903_o;
  wire [7:0] n10904_o;
  assign cy_o = n10903_o;
  assign ov_o = gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_n10893;
  assign rslt_o = n10904_o;
  /* addsub_core_struc.vhd:71:10  */
  assign s_cy = n10902_o; // (signal)
  /* addsub_core_struc.vhd:94:35  */
  assign n10879_o = opa_i[3:0];
  /* addsub_core_struc.vhd:95:35  */
  assign n10880_o = opb_i[3:0];
  /* addsub_core_struc.vhd:97:38  */
  assign n10881_o = s_cy[2];
  /* addsub_core_struc.vhd:98:29  */
  assign gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_n10882 = gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_cy_o; // (signal)
  /* addsub_core_struc.vhd:99:31  */
  assign gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_n10883 = gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_rslt_o; // (signal)
  /* addsub_core_struc.vhd:92:9  */
  addsub_cy_4 gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy (
    .opa_i(n10879_o),
    .opb_i(n10880_o),
    .addsub_i(addsub_i),
    .cy_i(n10881_o),
    .cy_o(gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_cy_o),
    .rslt_o(gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_rslt_o));
  /* addsub_core_struc.vhd:100:37  */
  assign n10888_o = s_cy[1];
  /* addsub_core_struc.vhd:105:35  */
  assign n10889_o = opa_i[7:4];
  /* addsub_core_struc.vhd:106:35  */
  assign n10890_o = opb_i[7:4];
  /* addsub_core_struc.vhd:108:49  */
  assign n10891_o = s_cy[1];
  /* addsub_core_struc.vhd:109:29  */
  assign gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_n10892 = gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_cy_o; // (signal)
  /* addsub_core_struc.vhd:110:29  */
  assign gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_n10893 = gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_ov_o; // (signal)
  /* addsub_core_struc.vhd:111:31  */
  assign gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_n10894 = gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_rslt_o; // (signal)
  /* addsub_core_struc.vhd:103:9  */
  addsub_ovcy_4 gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy (
    .opa_i(n10889_o),
    .opb_i(n10890_o),
    .addsub_i(addsub_i),
    .cy_i(n10891_o),
    .cy_o(gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_cy_o),
    .ov_o(gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_ov_o),
    .rslt_o(gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_rslt_o));
  assign n10902_o = {cy_i, gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_n10882, 1'bZ};
  assign n10903_o = {gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_n10892, n10888_o};
  assign n10904_o = {gen_greater_four_gen_addsub_n5_gen_last_addsub_i_addsub_ovcy_n10894, gen_greater_four_gen_addsub_n4_gen_nibble_addsub_i_addsub_cy_n10883};
endmodule

module alucore_8
  (input  [7:0] op_a_i,
   input  [7:0] op_b_i,
   input  [3:0] alu_cmd_i,
   input  [1:0] cy_i,
   output [1:0] cy_o,
   output [7:0] result_o);
  wire [7:0] n10784_o;
  wire n10786_o;
  wire [7:0] n10787_o;
  wire n10789_o;
  wire [7:0] n10790_o;
  wire n10792_o;
  wire [6:0] n10793_o;
  wire n10794_o;
  wire n10796_o;
  wire [6:0] n10797_o;
  wire n10798_o;
  wire n10799_o;
  wire n10800_o;
  wire n10802_o;
  wire [6:0] n10803_o;
  wire n10804_o;
  wire n10806_o;
  wire [6:0] n10807_o;
  wire n10808_o;
  wire n10809_o;
  wire n10810_o;
  wire n10812_o;
  wire n10813_o;
  wire [7:0] n10816_o;
  wire n10817_o;
  wire n10820_o;
  wire n10821_o;
  wire n10823_o;
  wire [7:0] n10824_o;
  wire n10826_o;
  wire [8:0] n10827_o;
  wire n10828_o;
  wire n10829_o;
  wire n10830_o;
  wire n10831_o;
  wire n10832_o;
  wire n10833_o;
  reg n10835_o;
  wire n10836_o;
  wire n10837_o;
  wire n10838_o;
  wire n10839_o;
  wire n10840_o;
  wire n10841_o;
  reg n10843_o;
  wire n10844_o;
  wire n10845_o;
  wire n10846_o;
  wire n10847_o;
  wire n10848_o;
  wire n10849_o;
  wire n10850_o;
  reg n10852_o;
  wire [5:0] n10853_o;
  wire [5:0] n10854_o;
  wire [5:0] n10855_o;
  wire [5:0] n10856_o;
  wire [5:0] n10857_o;
  wire [5:0] n10858_o;
  wire [5:0] n10859_o;
  wire [5:0] n10860_o;
  wire [5:0] n10861_o;
  reg [5:0] n10863_o;
  wire n10864_o;
  wire n10865_o;
  wire n10866_o;
  wire n10867_o;
  wire n10868_o;
  wire n10869_o;
  wire n10870_o;
  reg n10872_o;
  wire [1:0] n10874_o;
  wire [7:0] n10875_o;
  assign cy_o = n10874_o;
  assign result_o = n10875_o;
  /* alucore_rtl.vhd:86:26  */
  assign n10784_o = op_a_i & op_b_i;
  /* alucore_rtl.vhd:85:5  */
  assign n10786_o = alu_cmd_i == 4'b0011;
  /* alucore_rtl.vhd:90:26  */
  assign n10787_o = op_a_i | op_b_i;
  /* alucore_rtl.vhd:89:5  */
  assign n10789_o = alu_cmd_i == 4'b0101;
  /* alucore_rtl.vhd:94:26  */
  assign n10790_o = op_a_i ^ op_b_i;
  /* alucore_rtl.vhd:93:5  */
  assign n10792_o = alu_cmd_i == 4'b0110;
  /* alucore_rtl.vhd:99:46  */
  assign n10793_o = op_a_i[6:0];
  /* alucore_rtl.vhd:100:30  */
  assign n10794_o = op_a_i[7];
  /* alucore_rtl.vhd:97:5  */
  assign n10796_o = alu_cmd_i == 4'b0111;
  /* alucore_rtl.vhd:108:46  */
  assign n10797_o = op_a_i[6:0];
  /* alucore_rtl.vhd:109:28  */
  assign n10798_o = cy_i[1];
  /* alucore_rtl.vhd:114:35  */
  assign n10799_o = op_a_i[7];
  assign n10800_o = cy_i[0];
  /* alucore_rtl.vhd:106:5  */
  assign n10802_o = alu_cmd_i == 4'b1000;
  /* alucore_rtl.vhd:118:46  */
  assign n10803_o = op_a_i[7:1];
  /* alucore_rtl.vhd:119:37  */
  assign n10804_o = op_a_i[0];
  /* alucore_rtl.vhd:116:5  */
  assign n10806_o = alu_cmd_i == 4'b1001;
  /* alucore_rtl.vhd:127:46  */
  assign n10807_o = op_a_i[7:1];
  /* alucore_rtl.vhd:128:35  */
  assign n10808_o = cy_i[1];
  /* alucore_rtl.vhd:133:35  */
  assign n10809_o = op_a_i[0];
  assign n10810_o = cy_i[0];
  /* alucore_rtl.vhd:125:5  */
  assign n10812_o = alu_cmd_i == 4'b1010;
  /* alucore_rtl.vhd:136:17  */
  assign n10813_o = op_a_i == op_b_i;
  /* alucore_rtl.vhd:136:7  */
  assign n10816_o = n10813_o ? 8'b00000000 : 8'b11111111;
  /* alucore_rtl.vhd:142:17  */
  assign n10817_o = $unsigned(op_a_i) < $unsigned(op_b_i);
  /* alucore_rtl.vhd:142:7  */
  assign n10820_o = n10817_o ? 1'b1 : 1'b0;
  assign n10821_o = cy_i[0];
  /* alucore_rtl.vhd:135:5  */
  assign n10823_o = alu_cmd_i == 4'b1011;
  /* alucore_rtl.vhd:149:19  */
  assign n10824_o = ~op_a_i;
  /* alucore_rtl.vhd:148:5  */
  assign n10826_o = alu_cmd_i == 4'b1100;
  assign n10827_o = {n10826_o, n10823_o, n10812_o, n10806_o, n10802_o, n10796_o, n10792_o, n10789_o, n10786_o};
  assign n10828_o = cy_i[0];
  assign n10829_o = cy_i[0];
  assign n10830_o = cy_i[0];
  assign n10831_o = cy_i[0];
  assign n10832_o = cy_i[0];
  assign n10833_o = cy_i[0];
  /* alucore_rtl.vhd:83:3  */
  always @*
    case (n10827_o)
      9'b100000000: n10835_o = n10833_o;
      9'b010000000: n10835_o = n10821_o;
      9'b001000000: n10835_o = n10810_o;
      9'b000100000: n10835_o = n10832_o;
      9'b000010000: n10835_o = n10800_o;
      9'b000001000: n10835_o = n10831_o;
      9'b000000100: n10835_o = n10830_o;
      9'b000000010: n10835_o = n10829_o;
      9'b000000001: n10835_o = n10828_o;
      default: n10835_o = 1'b0;
    endcase
  assign n10836_o = cy_i[1];
  assign n10837_o = cy_i[1];
  assign n10838_o = cy_i[1];
  assign n10839_o = cy_i[1];
  assign n10840_o = cy_i[1];
  assign n10841_o = cy_i[1];
  /* alucore_rtl.vhd:83:3  */
  always @*
    case (n10827_o)
      9'b100000000: n10843_o = n10841_o;
      9'b010000000: n10843_o = n10820_o;
      9'b001000000: n10843_o = n10809_o;
      9'b000100000: n10843_o = n10840_o;
      9'b000010000: n10843_o = n10799_o;
      9'b000001000: n10843_o = n10839_o;
      9'b000000100: n10843_o = n10838_o;
      9'b000000010: n10843_o = n10837_o;
      9'b000000001: n10843_o = n10836_o;
      default: n10843_o = 1'b0;
    endcase
  assign n10844_o = n10784_o[0];
  assign n10845_o = n10787_o[0];
  assign n10846_o = n10790_o[0];
  assign n10847_o = n10803_o[0];
  assign n10848_o = n10807_o[0];
  assign n10849_o = n10816_o[0];
  assign n10850_o = n10824_o[0];
  /* alucore_rtl.vhd:83:3  */
  always @*
    case (n10827_o)
      9'b100000000: n10852_o = n10850_o;
      9'b010000000: n10852_o = n10849_o;
      9'b001000000: n10852_o = n10848_o;
      9'b000100000: n10852_o = n10847_o;
      9'b000010000: n10852_o = n10798_o;
      9'b000001000: n10852_o = n10794_o;
      9'b000000100: n10852_o = n10846_o;
      9'b000000010: n10852_o = n10845_o;
      9'b000000001: n10852_o = n10844_o;
      default: n10852_o = 1'b0;
    endcase
  assign n10853_o = n10784_o[6:1];
  assign n10854_o = n10787_o[6:1];
  assign n10855_o = n10790_o[6:1];
  assign n10856_o = n10793_o[5:0];
  assign n10857_o = n10797_o[5:0];
  assign n10858_o = n10803_o[6:1];
  assign n10859_o = n10807_o[6:1];
  assign n10860_o = n10816_o[6:1];
  assign n10861_o = n10824_o[6:1];
  /* alucore_rtl.vhd:83:3  */
  always @*
    case (n10827_o)
      9'b100000000: n10863_o = n10861_o;
      9'b010000000: n10863_o = n10860_o;
      9'b001000000: n10863_o = n10859_o;
      9'b000100000: n10863_o = n10858_o;
      9'b000010000: n10863_o = n10857_o;
      9'b000001000: n10863_o = n10856_o;
      9'b000000100: n10863_o = n10855_o;
      9'b000000010: n10863_o = n10854_o;
      9'b000000001: n10863_o = n10853_o;
      default: n10863_o = 6'b000000;
    endcase
  assign n10864_o = n10784_o[7];
  assign n10865_o = n10787_o[7];
  assign n10866_o = n10790_o[7];
  assign n10867_o = n10793_o[6];
  assign n10868_o = n10797_o[6];
  assign n10869_o = n10816_o[7];
  assign n10870_o = n10824_o[7];
  /* alucore_rtl.vhd:83:3  */
  always @*
    case (n10827_o)
      9'b100000000: n10872_o = n10870_o;
      9'b010000000: n10872_o = n10869_o;
      9'b001000000: n10872_o = n10808_o;
      9'b000100000: n10872_o = n10804_o;
      9'b000010000: n10872_o = n10868_o;
      9'b000001000: n10872_o = n10867_o;
      9'b000000100: n10872_o = n10866_o;
      9'b000000010: n10872_o = n10865_o;
      9'b000000001: n10872_o = n10864_o;
      default: n10872_o = 1'b0;
    endcase
  assign n10874_o = {n10843_o, n10835_o};
  assign n10875_o = {n10872_o, n10863_o, n10852_o};
endmodule

module alumux_8
  (input  [7:0] rom_data_i,
   input  [7:0] ram_data_i,
   input  [7:0] acc_i,
   input  [5:0] cmd_i,
   input  [1:0] cy_i,
   input  ov_i,
   input  [7:0] result_i,
   input  [1:0] new_cy_i,
   input  [7:0] addsub_rslt_i,
   input  [1:0] addsub_cy_i,
   input  addsub_ov_i,
   input  [7:0] qutnt_i,
   input  [7:0] rmndr_i,
   input  [15:0] product_i,
   input  [7:0] dcml_data_i,
   input  dcml_cy_i,
   output [1:0] cy_o,
   output ov_o,
   output [7:0] result_a_o,
   output [7:0] result_b_o,
   output [7:0] op_a_o,
   output [7:0] op_b_o,
   output [3:0] alu_cmd_o,
   output [7:0] opa_o,
   output [7:0] opb_o,
   output addsub_o,
   output addsub_cy_o,
   output [7:0] dvdnd_o,
   output [7:0] dvsor_o,
   output [7:0] mltplcnd_o,
   output [7:0] mltplctr_o,
   output [7:0] dcml_data_o);
  wire n10500_o;
  wire n10502_o;
  wire n10504_o;
  wire n10506_o;
  wire n10508_o;
  wire n10510_o;
  wire n10512_o;
  wire n10514_o;
  wire n10516_o;
  wire n10518_o;
  wire n10520_o;
  wire n10522_o;
  wire n10524_o;
  wire n10526_o;
  wire n10528_o;
  wire n10530_o;
  wire n10532_o;
  wire n10534_o;
  wire [17:0] n10535_o;
  reg [7:0] n10537_o;
  reg [7:0] n10545_o;
  reg [3:0] n10565_o;
  wire n10569_o;
  wire n10571_o;
  wire n10573_o;
  wire n10575_o;
  wire n10577_o;
  wire n10579_o;
  wire n10581_o;
  wire n10582_o;
  wire n10584_o;
  wire n10585_o;
  wire n10587_o;
  wire n10589_o;
  wire n10591_o;
  wire n10592_o;
  wire n10594_o;
  wire n10595_o;
  wire n10597_o;
  wire [12:0] n10598_o;
  reg [7:0] n10603_o;
  reg [7:0] n10612_o;
  reg n10627_o;
  reg n10638_o;
  reg [7:0] n10652_o;
  reg [7:0] n10666_o;
  reg [7:0] n10680_o;
  reg [7:0] n10694_o;
  reg [7:0] n10708_o;
  wire n10711_o;
  wire n10713_o;
  wire n10715_o;
  wire n10718_o;
  wire n10720_o;
  wire [7:0] n10721_o;
  wire [7:0] n10722_o;
  wire [7:0] n10723_o;
  wire n10725_o;
  wire n10728_o;
  wire n10730_o;
  wire n10732_o;
  wire n10734_o;
  wire n10735_o;
  wire n10737_o;
  wire n10738_o;
  wire n10740_o;
  wire n10741_o;
  wire n10743_o;
  wire n10744_o;
  wire n10746_o;
  wire n10747_o;
  wire n10749_o;
  wire n10751_o;
  wire n10752_o;
  wire n10754_o;
  wire n10755_o;
  wire n10757_o;
  wire n10758_o;
  wire [4:0] n10759_o;
  wire n10762_o;
  wire n10763_o;
  wire n10764_o;
  reg n10765_o;
  wire n10768_o;
  wire n10769_o;
  wire n10770_o;
  reg n10771_o;
  reg n10772_o;
  reg [7:0] n10773_o;
  reg [7:0] n10778_o;
  wire [1:0] n10780_o;
  assign cy_o = n10780_o;
  assign ov_o = n10772_o;
  assign result_a_o = n10773_o;
  assign result_b_o = n10778_o;
  assign op_a_o = n10537_o;
  assign op_b_o = n10545_o;
  assign alu_cmd_o = n10565_o;
  assign opa_o = n10603_o;
  assign opb_o = n10612_o;
  assign addsub_o = n10627_o;
  assign addsub_cy_o = n10638_o;
  assign dvdnd_o = n10652_o;
  assign dvsor_o = n10666_o;
  assign mltplcnd_o = n10680_o;
  assign mltplctr_o = n10694_o;
  assign dcml_data_o = n10708_o;
  /* alumux_rtl.vhd:119:8  */
  assign n10500_o = cmd_i == 6'b100101;
  /* alumux_rtl.vhd:123:8  */
  assign n10502_o = cmd_i == 6'b100110;
  /* alumux_rtl.vhd:127:8  */
  assign n10504_o = cmd_i == 6'b100111;
  /* alumux_rtl.vhd:131:8  */
  assign n10506_o = cmd_i == 6'b101100;
  /* alumux_rtl.vhd:135:8  */
  assign n10508_o = cmd_i == 6'b101101;
  /* alumux_rtl.vhd:139:8  */
  assign n10510_o = cmd_i == 6'b101110;
  /* alumux_rtl.vhd:143:8  */
  assign n10512_o = cmd_i == 6'b101111;
  /* alumux_rtl.vhd:147:8  */
  assign n10514_o = cmd_i == 6'b110000;
  /* alumux_rtl.vhd:151:8  */
  assign n10516_o = cmd_i == 6'b110001;
  /* alumux_rtl.vhd:155:8  */
  assign n10518_o = cmd_i == 6'b110010;
  /* alumux_rtl.vhd:159:8  */
  assign n10520_o = cmd_i == 6'b110011;
  /* alumux_rtl.vhd:163:8  */
  assign n10522_o = cmd_i == 6'b110100;
  /* alumux_rtl.vhd:167:8  */
  assign n10524_o = cmd_i == 6'b110101;
  /* alumux_rtl.vhd:171:8  */
  assign n10526_o = cmd_i == 6'b110110;
  /* alumux_rtl.vhd:175:8  */
  assign n10528_o = cmd_i == 6'b110111;
  /* alumux_rtl.vhd:179:8  */
  assign n10530_o = cmd_i == 6'b111010;
  /* alumux_rtl.vhd:183:8  */
  assign n10532_o = cmd_i == 6'b111011;
  /* alumux_rtl.vhd:187:8  */
  assign n10534_o = cmd_i == 6'b111100;
  assign n10535_o = {n10534_o, n10532_o, n10530_o, n10528_o, n10526_o, n10524_o, n10522_o, n10520_o, n10518_o, n10516_o, n10514_o, n10512_o, n10510_o, n10508_o, n10506_o, n10504_o, n10502_o, n10500_o};
  /* alumux_rtl.vhd:118:5  */
  always @*
    case (n10535_o)
      18'b100000000000000000: n10537_o = ram_data_i;
      18'b010000000000000000: n10537_o = acc_i;
      18'b001000000000000000: n10537_o = acc_i;
      18'b000100000000000000: n10537_o = ram_data_i;
      18'b000010000000000000: n10537_o = acc_i;
      18'b000001000000000000: n10537_o = acc_i;
      18'b000000100000000000: n10537_o = acc_i;
      18'b000000010000000000: n10537_o = acc_i;
      18'b000000001000000000: n10537_o = acc_i;
      18'b000000000100000000: n10537_o = rom_data_i;
      18'b000000000010000000: n10537_o = acc_i;
      18'b000000000001000000: n10537_o = acc_i;
      18'b000000000000100000: n10537_o = rom_data_i;
      18'b000000000000010000: n10537_o = acc_i;
      18'b000000000000001000: n10537_o = acc_i;
      18'b000000000000000100: n10537_o = ram_data_i;
      18'b000000000000000010: n10537_o = acc_i;
      18'b000000000000000001: n10537_o = acc_i;
      default: n10537_o = 8'b00000000;
    endcase
  /* alumux_rtl.vhd:118:5  */
  always @*
    case (n10535_o)
      18'b100000000000000000: n10545_o = rom_data_i;
      18'b010000000000000000: n10545_o = rom_data_i;
      18'b001000000000000000: n10545_o = ram_data_i;
      18'b000100000000000000: n10545_o = 8'b00000000;
      18'b000010000000000000: n10545_o = 8'b00000000;
      18'b000001000000000000: n10545_o = 8'b00000000;
      18'b000000100000000000: n10545_o = 8'b00000000;
      18'b000000010000000000: n10545_o = 8'b00000000;
      18'b000000001000000000: n10545_o = 8'b00000000;
      18'b000000000100000000: n10545_o = ram_data_i;
      18'b000000000010000000: n10545_o = rom_data_i;
      18'b000000000001000000: n10545_o = ram_data_i;
      18'b000000000000100000: n10545_o = ram_data_i;
      18'b000000000000010000: n10545_o = rom_data_i;
      18'b000000000000001000: n10545_o = ram_data_i;
      18'b000000000000000100: n10545_o = rom_data_i;
      18'b000000000000000010: n10545_o = rom_data_i;
      18'b000000000000000001: n10545_o = ram_data_i;
      default: n10545_o = 8'b00000000;
    endcase
  /* alumux_rtl.vhd:118:5  */
  always @*
    case (n10535_o)
      18'b100000000000000000: n10565_o = 4'b1011;
      18'b010000000000000000: n10565_o = 4'b1011;
      18'b001000000000000000: n10565_o = 4'b1011;
      18'b000100000000000000: n10565_o = 4'b1100;
      18'b000010000000000000: n10565_o = 4'b1100;
      18'b000001000000000000: n10565_o = 4'b1010;
      18'b000000100000000000: n10565_o = 4'b1001;
      18'b000000010000000000: n10565_o = 4'b1000;
      18'b000000001000000000: n10565_o = 4'b0111;
      18'b000000000100000000: n10565_o = 4'b0110;
      18'b000000000010000000: n10565_o = 4'b0110;
      18'b000000000001000000: n10565_o = 4'b0110;
      18'b000000000000100000: n10565_o = 4'b0101;
      18'b000000000000010000: n10565_o = 4'b0101;
      18'b000000000000001000: n10565_o = 4'b0101;
      18'b000000000000000100: n10565_o = 4'b0011;
      18'b000000000000000010: n10565_o = 4'b0011;
      18'b000000000000000001: n10565_o = 4'b0011;
      default: n10565_o = 4'b0000;
    endcase
  /* alumux_rtl.vhd:207:8  */
  assign n10569_o = cmd_i == 6'b100000;
  /* alumux_rtl.vhd:217:8  */
  assign n10571_o = cmd_i == 6'b101011;
  /* alumux_rtl.vhd:227:8  */
  assign n10573_o = cmd_i == 6'b101010;
  /* alumux_rtl.vhd:237:8  */
  assign n10575_o = cmd_i == 6'b111110;
  /* alumux_rtl.vhd:247:8  */
  assign n10577_o = cmd_i == 6'b111111;
  /* alumux_rtl.vhd:257:8  */
  assign n10579_o = cmd_i == 6'b111000;
  /* alumux_rtl.vhd:267:8  */
  assign n10581_o = cmd_i == 6'b111001;
  /* alumux_rtl.vhd:284:29  */
  assign n10582_o = cy_i[1];
  /* alumux_rtl.vhd:277:8  */
  assign n10584_o = cmd_i == 6'b101000;
  /* alumux_rtl.vhd:294:29  */
  assign n10585_o = cy_i[1];
  /* alumux_rtl.vhd:287:8  */
  assign n10587_o = cmd_i == 6'b101001;
  /* alumux_rtl.vhd:297:8  */
  assign n10589_o = cmd_i == 6'b100001;
  /* alumux_rtl.vhd:307:8  */
  assign n10591_o = cmd_i == 6'b100010;
  /* alumux_rtl.vhd:324:29  */
  assign n10592_o = cy_i[1];
  /* alumux_rtl.vhd:317:8  */
  assign n10594_o = cmd_i == 6'b100011;
  /* alumux_rtl.vhd:334:29  */
  assign n10595_o = cy_i[1];
  /* alumux_rtl.vhd:327:8  */
  assign n10597_o = cmd_i == 6'b100100;
  assign n10598_o = {n10597_o, n10594_o, n10591_o, n10589_o, n10587_o, n10584_o, n10581_o, n10579_o, n10577_o, n10575_o, n10573_o, n10571_o, n10569_o};
  /* alumux_rtl.vhd:206:5  */
  always @*
    case (n10598_o)
      13'b1000000000000: n10603_o = acc_i;
      13'b0100000000000: n10603_o = acc_i;
      13'b0010000000000: n10603_o = acc_i;
      13'b0001000000000: n10603_o = acc_i;
      13'b0000100000000: n10603_o = acc_i;
      13'b0000010000000: n10603_o = acc_i;
      13'b0000001000000: n10603_o = ram_data_i;
      13'b0000000100000: n10603_o = acc_i;
      13'b0000000010000: n10603_o = ram_data_i;
      13'b0000000001000: n10603_o = acc_i;
      13'b0000000000100: n10603_o = 8'b00000000;
      13'b0000000000010: n10603_o = 8'b00000000;
      13'b0000000000001: n10603_o = 8'b00000000;
      default: n10603_o = 8'b00000000;
    endcase
  /* alumux_rtl.vhd:206:5  */
  always @*
    case (n10598_o)
      13'b1000000000000: n10612_o = rom_data_i;
      13'b0100000000000: n10612_o = ram_data_i;
      13'b0010000000000: n10612_o = rom_data_i;
      13'b0001000000000: n10612_o = ram_data_i;
      13'b0000100000000: n10612_o = rom_data_i;
      13'b0000010000000: n10612_o = ram_data_i;
      13'b0000001000000: n10612_o = 8'b00000001;
      13'b0000000100000: n10612_o = 8'b00000001;
      13'b0000000010000: n10612_o = 8'b00000001;
      13'b0000000001000: n10612_o = 8'b00000001;
      13'b0000000000100: n10612_o = 8'b00000000;
      13'b0000000000010: n10612_o = 8'b00000000;
      13'b0000000000001: n10612_o = 8'b00000000;
      default: n10612_o = 8'b00000000;
    endcase
  /* alumux_rtl.vhd:206:5  */
  always @*
    case (n10598_o)
      13'b1000000000000: n10627_o = 1'b1;
      13'b0100000000000: n10627_o = 1'b1;
      13'b0010000000000: n10627_o = 1'b1;
      13'b0001000000000: n10627_o = 1'b1;
      13'b0000100000000: n10627_o = 1'b0;
      13'b0000010000000: n10627_o = 1'b0;
      13'b0000001000000: n10627_o = 1'b0;
      13'b0000000100000: n10627_o = 1'b0;
      13'b0000000010000: n10627_o = 1'b1;
      13'b0000000001000: n10627_o = 1'b1;
      13'b0000000000100: n10627_o = 1'b0;
      13'b0000000000010: n10627_o = 1'b0;
      13'b0000000000001: n10627_o = 1'b0;
      default: n10627_o = 1'b0;
    endcase
  /* alumux_rtl.vhd:206:5  */
  always @*
    case (n10598_o)
      13'b1000000000000: n10638_o = n10595_o;
      13'b0100000000000: n10638_o = n10592_o;
      13'b0010000000000: n10638_o = 1'b0;
      13'b0001000000000: n10638_o = 1'b0;
      13'b0000100000000: n10638_o = n10585_o;
      13'b0000010000000: n10638_o = n10582_o;
      13'b0000001000000: n10638_o = 1'b0;
      13'b0000000100000: n10638_o = 1'b0;
      13'b0000000010000: n10638_o = 1'b0;
      13'b0000000001000: n10638_o = 1'b0;
      13'b0000000000100: n10638_o = 1'b0;
      13'b0000000000010: n10638_o = 1'b0;
      13'b0000000000001: n10638_o = 1'b0;
      default: n10638_o = 1'b0;
    endcase
  /* alumux_rtl.vhd:206:5  */
  always @*
    case (n10598_o)
      13'b1000000000000: n10652_o = 8'b00000000;
      13'b0100000000000: n10652_o = 8'b00000000;
      13'b0010000000000: n10652_o = 8'b00000000;
      13'b0001000000000: n10652_o = 8'b00000000;
      13'b0000100000000: n10652_o = 8'b00000000;
      13'b0000010000000: n10652_o = 8'b00000000;
      13'b0000001000000: n10652_o = 8'b00000000;
      13'b0000000100000: n10652_o = 8'b00000000;
      13'b0000000010000: n10652_o = 8'b00000000;
      13'b0000000001000: n10652_o = 8'b00000000;
      13'b0000000000100: n10652_o = 8'b00000000;
      13'b0000000000010: n10652_o = acc_i;
      13'b0000000000001: n10652_o = 8'b00000000;
      default: n10652_o = 8'b00000000;
    endcase
  /* alumux_rtl.vhd:206:5  */
  always @*
    case (n10598_o)
      13'b1000000000000: n10666_o = 8'b00000000;
      13'b0100000000000: n10666_o = 8'b00000000;
      13'b0010000000000: n10666_o = 8'b00000000;
      13'b0001000000000: n10666_o = 8'b00000000;
      13'b0000100000000: n10666_o = 8'b00000000;
      13'b0000010000000: n10666_o = 8'b00000000;
      13'b0000001000000: n10666_o = 8'b00000000;
      13'b0000000100000: n10666_o = 8'b00000000;
      13'b0000000010000: n10666_o = 8'b00000000;
      13'b0000000001000: n10666_o = 8'b00000000;
      13'b0000000000100: n10666_o = 8'b00000000;
      13'b0000000000010: n10666_o = ram_data_i;
      13'b0000000000001: n10666_o = 8'b00000000;
      default: n10666_o = 8'b00000000;
    endcase
  /* alumux_rtl.vhd:206:5  */
  always @*
    case (n10598_o)
      13'b1000000000000: n10680_o = 8'b00000000;
      13'b0100000000000: n10680_o = 8'b00000000;
      13'b0010000000000: n10680_o = 8'b00000000;
      13'b0001000000000: n10680_o = 8'b00000000;
      13'b0000100000000: n10680_o = 8'b00000000;
      13'b0000010000000: n10680_o = 8'b00000000;
      13'b0000001000000: n10680_o = 8'b00000000;
      13'b0000000100000: n10680_o = 8'b00000000;
      13'b0000000010000: n10680_o = 8'b00000000;
      13'b0000000001000: n10680_o = 8'b00000000;
      13'b0000000000100: n10680_o = acc_i;
      13'b0000000000010: n10680_o = 8'b00000000;
      13'b0000000000001: n10680_o = 8'b00000000;
      default: n10680_o = 8'b00000000;
    endcase
  /* alumux_rtl.vhd:206:5  */
  always @*
    case (n10598_o)
      13'b1000000000000: n10694_o = 8'b00000000;
      13'b0100000000000: n10694_o = 8'b00000000;
      13'b0010000000000: n10694_o = 8'b00000000;
      13'b0001000000000: n10694_o = 8'b00000000;
      13'b0000100000000: n10694_o = 8'b00000000;
      13'b0000010000000: n10694_o = 8'b00000000;
      13'b0000001000000: n10694_o = 8'b00000000;
      13'b0000000100000: n10694_o = 8'b00000000;
      13'b0000000010000: n10694_o = 8'b00000000;
      13'b0000000001000: n10694_o = 8'b00000000;
      13'b0000000000100: n10694_o = ram_data_i;
      13'b0000000000010: n10694_o = 8'b00000000;
      13'b0000000000001: n10694_o = 8'b00000000;
      default: n10694_o = 8'b00000000;
    endcase
  /* alumux_rtl.vhd:206:5  */
  always @*
    case (n10598_o)
      13'b1000000000000: n10708_o = 8'b00000000;
      13'b0100000000000: n10708_o = 8'b00000000;
      13'b0010000000000: n10708_o = 8'b00000000;
      13'b0001000000000: n10708_o = 8'b00000000;
      13'b0000100000000: n10708_o = 8'b00000000;
      13'b0000010000000: n10708_o = 8'b00000000;
      13'b0000001000000: n10708_o = 8'b00000000;
      13'b0000000100000: n10708_o = 8'b00000000;
      13'b0000000010000: n10708_o = 8'b00000000;
      13'b0000000001000: n10708_o = 8'b00000000;
      13'b0000000000100: n10708_o = 8'b00000000;
      13'b0000000000010: n10708_o = 8'b00000000;
      13'b0000000000001: n10708_o = acc_i;
      default: n10708_o = 8'b00000000;
    endcase
  assign n10711_o = cy_i[0];
  /* alumux_rtl.vhd:367:8  */
  assign n10713_o = cmd_i == 6'b100000;
  /* alumux_rtl.vhd:385:26  */
  assign n10715_o = ram_data_i == 8'b00000000;
  /* alumux_rtl.vhd:385:12  */
  assign n10718_o = n10715_o ? 1'b1 : 1'b0;
  /* alumux_rtl.vhd:380:8  */
  assign n10720_o = cmd_i == 6'b101011;
  /* alumux_rtl.vhd:398:43  */
  assign n10721_o = product_i[7:0];
  /* alumux_rtl.vhd:399:43  */
  assign n10722_o = product_i[15:8];
  /* alumux_rtl.vhd:401:24  */
  assign n10723_o = product_i[15:8];
  /* alumux_rtl.vhd:402:16  */
  assign n10725_o = n10723_o == 8'b00000000;
  /* alumux_rtl.vhd:401:12  */
  assign n10728_o = n10725_o ? 1'b0 : 1'b1;
  /* alumux_rtl.vhd:396:8  */
  assign n10730_o = cmd_i == 6'b101010;
  /* alumux_rtl.vhd:413:8  */
  assign n10732_o = cmd_i == 6'b101000;
  /* alumux_rtl.vhd:413:25  */
  assign n10734_o = cmd_i == 6'b101001;
  /* alumux_rtl.vhd:413:25  */
  assign n10735_o = n10732_o | n10734_o;
  /* alumux_rtl.vhd:413:39  */
  assign n10737_o = cmd_i == 6'b100001;
  /* alumux_rtl.vhd:413:39  */
  assign n10738_o = n10735_o | n10737_o;
  /* alumux_rtl.vhd:413:53  */
  assign n10740_o = cmd_i == 6'b100010;
  /* alumux_rtl.vhd:413:53  */
  assign n10741_o = n10738_o | n10740_o;
  /* alumux_rtl.vhd:413:67  */
  assign n10743_o = cmd_i == 6'b100011;
  /* alumux_rtl.vhd:413:67  */
  assign n10744_o = n10741_o | n10743_o;
  /* alumux_rtl.vhd:414:26  */
  assign n10746_o = cmd_i == 6'b100100;
  /* alumux_rtl.vhd:414:26  */
  assign n10747_o = n10744_o | n10746_o;
  /* alumux_rtl.vhd:419:8  */
  assign n10749_o = cmd_i == 6'b111110;
  /* alumux_rtl.vhd:419:21  */
  assign n10751_o = cmd_i == 6'b111111;
  /* alumux_rtl.vhd:419:21  */
  assign n10752_o = n10749_o | n10751_o;
  /* alumux_rtl.vhd:419:31  */
  assign n10754_o = cmd_i == 6'b111000;
  /* alumux_rtl.vhd:419:31  */
  assign n10755_o = n10752_o | n10754_o;
  /* alumux_rtl.vhd:419:41  */
  assign n10757_o = cmd_i == 6'b111001;
  /* alumux_rtl.vhd:419:41  */
  assign n10758_o = n10755_o | n10757_o;
  assign n10759_o = {n10758_o, n10747_o, n10730_o, n10720_o, n10713_o};
  assign n10762_o = addsub_cy_i[0];
  assign n10763_o = cy_i[0];
  assign n10764_o = new_cy_i[0];
  /* alumux_rtl.vhd:366:5  */
  always @*
    case (n10759_o)
      5'b10000: n10765_o = n10763_o;
      5'b01000: n10765_o = n10762_o;
      5'b00100: n10765_o = 1'b0;
      5'b00010: n10765_o = 1'b0;
      5'b00001: n10765_o = n10711_o;
      default: n10765_o = n10764_o;
    endcase
  assign n10768_o = addsub_cy_i[1];
  assign n10769_o = cy_i[1];
  assign n10770_o = new_cy_i[1];
  /* alumux_rtl.vhd:366:5  */
  always @*
    case (n10759_o)
      5'b10000: n10771_o = n10769_o;
      5'b01000: n10771_o = n10768_o;
      5'b00100: n10771_o = 1'b0;
      5'b00010: n10771_o = 1'b0;
      5'b00001: n10771_o = dcml_cy_i;
      default: n10771_o = n10770_o;
    endcase
  /* alumux_rtl.vhd:366:5  */
  always @*
    case (n10759_o)
      5'b10000: n10772_o = addsub_ov_i;
      5'b01000: n10772_o = addsub_ov_i;
      5'b00100: n10772_o = n10728_o;
      5'b00010: n10772_o = n10718_o;
      5'b00001: n10772_o = ov_i;
      default: n10772_o = ov_i;
    endcase
  /* alumux_rtl.vhd:366:5  */
  always @*
    case (n10759_o)
      5'b10000: n10773_o = addsub_rslt_i;
      5'b01000: n10773_o = addsub_rslt_i;
      5'b00100: n10773_o = n10721_o;
      5'b00010: n10773_o = qutnt_i;
      5'b00001: n10773_o = dcml_data_i;
      default: n10773_o = result_i;
    endcase
  /* alumux_rtl.vhd:366:5  */
  always @*
    case (n10759_o)
      5'b10000: n10778_o = 8'b00000000;
      5'b01000: n10778_o = 8'b00000000;
      5'b00100: n10778_o = n10722_o;
      5'b00010: n10778_o = rmndr_i;
      5'b00001: n10778_o = 8'b00000000;
      default: n10778_o = 8'b00000000;
    endcase
  assign n10780_o = {n10771_o, n10765_o};
endmodule

module control_mem
  (input  [7:0] rom_data_i,
   input  [7:0] ram_data_i,
   input  [7:0] aludata_i,
   input  [7:0] aludatb_i,
   input  [1:0] new_cy_i,
   input  new_ov_i,
   input  reset,
   input  clk,
   input  cen,
   input  int0_i,
   input  int1_i,
   input  [7:0] p0_i,
   input  [7:0] p1_i,
   input  [7:0] p2_i,
   input  [7:0] p3_i,
   input  [2:0] all_scon_i,
   input  [7:0] all_sbuf_i,
   input  all_tf0_i,
   input  all_tf1_i,
   input  [7:0] all_tl0_i,
   input  [7:0] all_tl1_i,
   input  [7:0] all_th0_i,
   input  [7:0] all_th1_i,
   input  [7:0] datax_i,
   input  [3:0] pc_inc_en_i,
   input  [2:0] nextstate_i,
   input  [3:0] adr_mux_i,
   input  [1:0] adrx_mux_i,
   input  wrx_mux_i,
   input  [3:0] data_mux_i,
   input  [3:0] bdata_mux_i,
   input  [2:0] regs_wr_en_i,
   input  [3:0] help_en_i,
   input  [1:0] help16_en_i,
   input  helpb_en_i,
   input  inthigh_en_i,
   input  intlow_en_i,
   input  intpre2_en_i,
   input  inthigh_d_i,
   input  intlow_d_i,
   input  intpre2_d_i,
   input  ext0isr_d_i,
   input  ext1isr_d_i,
   input  ext0isrh_d_i,
   input  ext1isrh_d_i,
   input  ext0isr_en_i,
   input  ext1isr_en_i,
   input  ext0isrh_en_i,
   input  ext1isrh_en_i,
   output [15:0] pc_o,
   output [7:0] ram_data_o,
   output [6:0] ram_adr_o,
   output [7:0] reg_data_o,
   output ram_wr_o,
   output [1:0] cy_o,
   output ov_o,
   output ram_en_o,
   output [7:0] acc_o,
   output [7:0] p0_o,
   output [7:0] p1_o,
   output [7:0] p2_o,
   output [7:0] p3_o,
   output all_trans_o,
   output [5:0] all_scon_o,
   output [7:0] all_sbuf_o,
   output all_smod_o,
   output all_tcon_tr0_o,
   output all_tcon_tr1_o,
   output [7:0] all_tmod_o,
   output [7:0] all_reload_o,
   output [1:0] all_wt_o,
   output all_wt_en_o,
   output [2:0] state_o,
   output [7:0] help_o,
   output bit_data_o,
   output [7:0] command_o,
   output inthigh_o,
   output intlow_o,
   output intpre_o,
   output intpre2_o,
   output intblock_o,
   output ti_o,
   output ri_o,
   output ie0_o,
   output ie1_o,
   output tf0_o,
   output tf1_o,
   output [7:0] psw_o,
   output [7:0] ie_o,
   output [7:0] ip_o,
   output [15:0] adrx_o,
   output [7:0] datax_o,
   output wrx_o,
   output memx_o);
  wire [7:0] s_help;
  wire [15:0] s_help16;
  wire s_helpb;
  wire [7:0] s_ir;
  wire [127:0] gprbit;
  wire [7:0] s_r0_b0;
  wire [7:0] s_r1_b0;
  wire [7:0] s_r0_b1;
  wire [7:0] s_r1_b1;
  wire [7:0] s_r0_b2;
  wire [7:0] s_r1_b2;
  wire [7:0] s_r0_b3;
  wire [7:0] s_r1_b3;
  wire [7:0] s_reg_data;
  wire [2:0] state;
  wire [7:0] s_command;
  wire [3:0] s_pc_inc_en;
  wire [2:0] s_regs_wr_en;
  wire [3:0] s_data_mux;
  wire [3:0] s_bdata_mux;
  wire [3:0] s_adr_mux;
  wire [1:0] s_adrx_mux;
  wire [3:0] s_help_en;
  wire [1:0] s_help16_en;
  wire s_helpb_en;
  wire s_intpre2_d;
  wire s_intpre2_en;
  wire s_intlow_d;
  wire s_intlow_en;
  wire s_inthigh_d;
  wire s_inthigh_en;
  wire s_ext0isr_d;
  wire s_ext0isrh_d;
  wire s_ext1isr_d;
  wire s_ext1isrh_d;
  wire [2:0] s_nextstate;
  wire s_bit_data;
  wire s_intpre;
  wire s_intpre2;
  wire s_inthigh;
  wire s_intlow;
  wire s_intblock;
  wire s_intblock_o;
  wire s_int0_edge;
  wire s_int1_edge;
  wire s_tf0_edge;
  wire s_tf1_edge;
  wire s_ri_edge;
  wire s_ti_edge;
  wire s_smodreg;
  wire [7:0] s_tl0;
  wire [7:0] s_tl1;
  wire [7:0] s_th0;
  wire [7:0] s_th1;
  wire [7:0] s_sbufi;
  wire [7:0] s_reload;
  wire [1:0] s_wt;
  wire s_tf1;
  wire s_tf0;
  wire s_ie1;
  wire s_ie0;
  wire s_ri;
  wire s_ti;
  wire s_rb8;
  wire s_tb8;
  wire s_ren;
  wire s_sm2;
  wire s_sm1;
  wire s_sm0;
  wire s_smod;
  wire s_int0_h1;
  wire s_int0_h2;
  wire s_int0_h3;
  wire s_int1_h1;
  wire s_int1_h2;
  wire s_int1_h3;
  wire s_tf0_h1;
  wire s_tf0_h2;
  wire s_tf1_h1;
  wire s_tf1_h2;
  wire s_ri_h1;
  wire s_ri_h2;
  wire s_ti_h1;
  wire s_ti_h2;
  wire s_p;
  wire [7:0] s_p0;
  wire [7:0] s_p1;
  wire [7:0] s_p2;
  wire [7:0] s_p3;
  wire [15:0] pc;
  wire [15:0] pc_comb;
  wire [15:0] pc_plus1;
  wire [15:0] pc_plus2;
  wire [7:0] s_data;
  wire [7:0] s_adr;
  wire [7:0] s_preadr;
  wire s_bdata;
  wire [7:0] s_rr_adr;
  wire [7:0] s_ri_adr;
  wire [7:0] s_ri_data;
  wire [7:0] p0;
  wire [7:0] sp;
  wire [7:0] dpl;
  wire [7:0] dph;
  wire [3:0] pcon;
  wire [7:0] tcon;
  wire [7:0] tmod;
  wire [7:0] p1;
  wire [7:0] scon;
  wire [7:0] sbuf;
  wire [7:0] p2;
  wire [7:0] ie;
  wire [7:0] p3;
  wire [7:0] ip;
  wire [7:0] psw;
  wire [7:0] acc;
  wire [7:0] b;
  wire [7:0] tsel;
  wire [7:0] ssel;
  wire [15:0] n7280_o;
  wire [15:0] n7283_o;
  wire [6:0] n7284_o;
  wire n7285_o;
  wire n7286_o;
  wire n7287_o;
  wire n7302_o;
  wire n7303_o;
  wire n7304_o;
  wire n7305_o;
  wire n7306_o;
  wire n7307_o;
  wire n7308_o;
  wire n7309_o;
  wire n7310_o;
  wire n7311_o;
  wire n7312_o;
  wire n7313_o;
  wire n7314_o;
  wire n7315_o;
  wire n7316_o;
  wire n7317_o;
  wire n7318_o;
  wire n7319_o;
  wire n7320_o;
  wire n7321_o;
  wire n7322_o;
  wire n7323_o;
  wire n7324_o;
  wire n7325_o;
  wire n7326_o;
  wire n7327_o;
  wire n7328_o;
  wire n7329_o;
  wire n7330_o;
  wire n7331_o;
  wire n7332_o;
  wire n7333_o;
  wire n7334_o;
  wire n7335_o;
  wire n7336_o;
  wire n7338_o;
  wire [7:0] n7339_o;
  wire [7:0] n7341_o;
  wire [7:0] n7343_o;
  wire [7:0] n7344_o;
  wire [7:0] n7346_o;
  wire [7:0] n7348_o;
  wire [7:0] n7349_o;
  wire n7353_o;
  wire n7355_o;
  wire [31:0] n7356_o;
  wire n7358_o;
  wire [31:0] n7359_o;
  wire n7361_o;
  wire n7362_o;
  wire n7363_o;
  wire n7364_o;
  wire n7365_o;
  wire n7366_o;
  wire n7368_o;
  wire [4:0] n7369_o;
  wire n7371_o;
  wire [4:0] n7372_o;
  wire n7374_o;
  wire n7375_o;
  wire n7376_o;
  wire n7377_o;
  wire n7378_o;
  wire n7379_o;
  wire n7381_o;
  wire n7383_o;
  wire n7384_o;
  wire n7386_o;
  wire n7388_o;
  wire n7391_o;
  wire [31:0] n7392_o;
  wire n7394_o;
  wire n7396_o;
  wire n7398_o;
  wire n7400_o;
  localparam [2:0] n7401_o = 3'b000;
  wire n7403_o;
  wire n7405_o;
  wire n7407_o;
  wire n7409_o;
  wire n7411_o;
  wire n7413_o;
  wire n7415_o;
  wire n7417_o;
  wire n7419_o;
  wire n7421_o;
  wire n7423_o;
  wire n7425_o;
  wire n7427_o;
  wire n7429_o;
  wire n7431_o;
  wire n7433_o;
  wire n7435_o;
  wire n7437_o;
  wire n7439_o;
  wire [22:0] n7440_o;
  wire n7441_o;
  wire n7442_o;
  wire n7443_o;
  wire n7444_o;
  wire n7445_o;
  wire n7446_o;
  wire n7447_o;
  wire n7448_o;
  wire n7449_o;
  wire n7450_o;
  wire n7451_o;
  wire n7452_o;
  wire n7453_o;
  wire n7454_o;
  wire n7455_o;
  wire n7456_o;
  wire n7457_o;
  wire n7458_o;
  wire n7459_o;
  wire n7460_o;
  wire n7461_o;
  wire n7462_o;
  reg n7464_o;
  wire n7465_o;
  wire n7466_o;
  wire n7467_o;
  wire n7468_o;
  wire n7469_o;
  wire n7470_o;
  wire n7471_o;
  wire n7472_o;
  wire n7473_o;
  wire n7474_o;
  wire n7475_o;
  wire n7476_o;
  wire n7477_o;
  wire n7478_o;
  wire n7479_o;
  wire n7480_o;
  wire n7481_o;
  wire n7482_o;
  wire n7483_o;
  wire n7484_o;
  wire n7485_o;
  wire n7486_o;
  reg n7488_o;
  wire n7489_o;
  wire n7490_o;
  wire n7491_o;
  wire n7492_o;
  wire n7493_o;
  wire n7494_o;
  wire n7495_o;
  wire n7496_o;
  wire n7497_o;
  wire n7498_o;
  wire n7499_o;
  wire n7500_o;
  wire n7501_o;
  wire n7502_o;
  wire n7503_o;
  wire n7504_o;
  wire n7505_o;
  wire n7506_o;
  wire n7507_o;
  wire n7508_o;
  wire n7509_o;
  wire n7510_o;
  reg n7512_o;
  wire n7513_o;
  wire n7514_o;
  wire n7515_o;
  wire n7516_o;
  wire n7517_o;
  wire n7518_o;
  wire n7519_o;
  wire n7520_o;
  wire n7521_o;
  wire n7522_o;
  wire n7523_o;
  wire n7524_o;
  wire n7525_o;
  wire n7526_o;
  wire n7527_o;
  wire n7528_o;
  wire n7529_o;
  wire n7530_o;
  wire n7531_o;
  wire n7532_o;
  wire n7533_o;
  wire n7534_o;
  reg n7536_o;
  wire n7537_o;
  wire n7538_o;
  wire n7539_o;
  wire n7540_o;
  wire n7541_o;
  wire n7542_o;
  wire n7543_o;
  wire n7544_o;
  wire n7545_o;
  wire n7546_o;
  wire n7547_o;
  wire n7548_o;
  wire n7549_o;
  wire n7550_o;
  wire n7551_o;
  wire n7552_o;
  wire n7553_o;
  wire n7554_o;
  wire n7555_o;
  wire n7556_o;
  wire n7557_o;
  wire n7558_o;
  reg n7560_o;
  wire n7561_o;
  wire n7562_o;
  wire n7563_o;
  wire n7564_o;
  wire n7565_o;
  wire n7566_o;
  wire n7567_o;
  wire n7568_o;
  wire n7569_o;
  wire n7570_o;
  wire n7571_o;
  wire n7572_o;
  wire n7573_o;
  wire n7574_o;
  wire n7575_o;
  wire n7576_o;
  wire n7577_o;
  wire n7578_o;
  wire n7579_o;
  wire n7580_o;
  wire n7581_o;
  wire n7582_o;
  reg n7584_o;
  wire n7585_o;
  wire n7586_o;
  wire n7587_o;
  wire n7588_o;
  wire n7589_o;
  wire n7590_o;
  wire n7591_o;
  wire n7592_o;
  wire n7593_o;
  wire n7594_o;
  wire n7595_o;
  wire n7596_o;
  wire n7597_o;
  wire n7598_o;
  wire n7599_o;
  wire n7600_o;
  wire n7601_o;
  wire n7602_o;
  wire n7603_o;
  wire n7604_o;
  wire n7605_o;
  wire n7606_o;
  reg n7608_o;
  wire n7609_o;
  wire n7610_o;
  wire n7611_o;
  wire n7612_o;
  wire n7613_o;
  wire n7614_o;
  wire n7615_o;
  wire n7616_o;
  wire n7617_o;
  wire n7618_o;
  wire n7619_o;
  wire n7620_o;
  wire n7621_o;
  wire n7622_o;
  wire n7623_o;
  wire n7624_o;
  wire n7625_o;
  wire n7626_o;
  wire n7627_o;
  wire n7628_o;
  wire n7629_o;
  reg n7631_o;
  wire [3:0] n7632_o;
  wire n7634_o;
  wire [3:0] n7635_o;
  wire n7640_o;
  wire n7642_o;
  wire n7644_o;
  wire n7646_o;
  wire n7648_o;
  wire n7650_o;
  wire n7652_o;
  wire n7654_o;
  wire [7:0] n7655_o;
  wire [7:0] n7656_o;
  wire [7:0] n7657_o;
  wire [7:0] n7658_o;
  wire [7:0] n7659_o;
  wire [7:0] n7660_o;
  wire [7:0] n7661_o;
  wire [7:0] n7662_o;
  wire [7:0] n7663_o;
  wire [7:0] n7664_o;
  wire [7:0] n7665_o;
  wire n7666_o;
  wire [3:0] n7667_o;
  wire [2:0] n7668_o;
  wire n7673_o;
  wire [2:0] n7674_o;
  wire n7679_o;
  wire [2:0] n7680_o;
  wire n7685_o;
  wire [2:0] n7686_o;
  wire [31:0] n7687_o;
  wire n7689_o;
  wire [2:0] n7690_o;
  wire n7694_o;
  wire n7696_o;
  wire [2:0] n7697_o;
  wire n7702_o;
  wire [2:0] n7703_o;
  wire n7708_o;
  wire [2:0] n7709_o;
  wire n7714_o;
  wire [2:0] n7715_o;
  wire n7720_o;
  wire [2:0] n7721_o;
  wire n7726_o;
  wire [2:0] n7727_o;
  wire n7732_o;
  wire [2:0] n7733_o;
  wire n7738_o;
  wire [10:0] n7739_o;
  reg n7741_o;
  wire [3:0] n7742_o;
  wire [2:0] n7745_o;
  wire n7750_o;
  wire n7752_o;
  wire n7753_o;
  wire n7754_o;
  wire n7755_o;
  wire n7756_o;
  wire n7757_o;
  wire n7758_o;
  wire n7759_o;
  wire n7760_o;
  wire n7761_o;
  wire n7762_o;
  wire n7763_o;
  wire n7767_o;
  wire n7768_o;
  wire n7816_o;
  wire n7817_o;
  wire n7818_o;
  wire n7819_o;
  wire n7820_o;
  wire n7821_o;
  wire n7822_o;
  wire n7823_o;
  wire n7824_o;
  wire n7825_o;
  wire n7826_o;
  wire n7827_o;
  wire n7828_o;
  wire n7829_o;
  wire n7830_o;
  wire n7831_o;
  wire n7832_o;
  wire n7833_o;
  wire n7834_o;
  wire n7835_o;
  wire n7836_o;
  wire n7837_o;
  wire n7838_o;
  wire n7839_o;
  wire n7840_o;
  wire n7841_o;
  wire n7842_o;
  wire n7843_o;
  wire n7844_o;
  wire n7845_o;
  wire n7846_o;
  wire n7847_o;
  wire n7848_o;
  wire n7849_o;
  wire n7850_o;
  wire n7851_o;
  wire n7854_o;
  wire n7855_o;
  wire n7856_o;
  wire n7857_o;
  wire n7858_o;
  wire n7859_o;
  wire n7860_o;
  wire n7861_o;
  wire n7862_o;
  wire n7863_o;
  wire n7864_o;
  wire n7865_o;
  wire n7866_o;
  wire n7867_o;
  wire n7868_o;
  wire n7869_o;
  wire n7872_o;
  wire n7873_o;
  wire n7875_o;
  wire n7877_o;
  wire n7881_o;
  wire [7:0] n7882_o;
  wire n7884_o;
  wire [7:0] n7885_o;
  wire n7887_o;
  wire n7889_o;
  wire n7891_o;
  wire n7893_o;
  wire n7895_o;
  wire [3:0] n7896_o;
  wire [3:0] n7897_o;
  wire n7899_o;
  wire n7901_o;
  wire [3:0] n7902_o;
  wire [3:0] n7903_o;
  wire n7905_o;
  wire [3:0] n7906_o;
  wire [3:0] n7907_o;
  wire n7909_o;
  wire [7:0] n7910_o;
  wire n7912_o;
  wire [7:0] n7913_o;
  wire n7915_o;
  wire [7:0] n7916_o;
  wire n7918_o;
  wire n7920_o;
  wire [14:0] n7921_o;
  wire [3:0] n7923_o;
  wire [3:0] n7924_o;
  wire [3:0] n7925_o;
  wire [3:0] n7926_o;
  wire [3:0] n7927_o;
  wire [3:0] n7928_o;
  wire [3:0] n7929_o;
  wire [3:0] n7930_o;
  wire [3:0] n7931_o;
  wire [3:0] n7932_o;
  wire [3:0] n7933_o;
  reg [3:0] n7935_o;
  wire [3:0] n7937_o;
  wire [3:0] n7938_o;
  wire [3:0] n7939_o;
  wire [3:0] n7940_o;
  wire [3:0] n7941_o;
  wire [3:0] n7942_o;
  wire [3:0] n7943_o;
  wire [3:0] n7944_o;
  wire [3:0] n7945_o;
  wire [3:0] n7946_o;
  wire [3:0] n7947_o;
  reg [3:0] n7949_o;
  wire n7951_o;
  wire n7952_o;
  wire n7953_o;
  wire n7955_o;
  wire n7956_o;
  wire n7957_o;
  wire n7958_o;
  wire n7960_o;
  wire n7961_o;
  wire n7963_o;
  wire n7965_o;
  wire n7966_o;
  wire n7967_o;
  wire n7969_o;
  wire n7970_o;
  wire n7972_o;
  wire n7974_o;
  wire n7975_o;
  wire n7977_o;
  wire n7978_o;
  wire n7979_o;
  wire n7981_o;
  wire n7982_o;
  wire n7983_o;
  wire n7984_o;
  wire n7986_o;
  wire n7988_o;
  wire [11:0] n7989_o;
  reg n7993_o;
  wire n7995_o;
  wire n7997_o;
  wire n7999_o;
  wire n8001_o;
  wire n8003_o;
  wire n8005_o;
  wire n8007_o;
  wire n8009_o;
  wire n8011_o;
  wire n8013_o;
  wire n8015_o;
  wire n8017_o;
  wire n8019_o;
  wire n8021_o;
  wire n8023_o;
  wire [7:0] n8026_o;
  wire n8028_o;
  wire [15:0] n8029_o;
  reg [7:0] n8040_o;
  wire n8042_o;
  wire n8045_o;
  wire [1:0] n8046_o;
  reg [7:0] n8048_o;
  reg [7:0] n8050_o;
  reg n8054_o;
  wire n8056_o;
  wire n8058_o;
  wire n8060_o;
  wire n8062_o;
  wire n8064_o;
  wire n8066_o;
  wire n8068_o;
  wire n8070_o;
  wire [7:0] n8071_o;
  reg [7:0] n8073_o;
  wire n8075_o;
  wire n8077_o;
  wire n8078_o;
  wire n8079_o;
  wire [3:0] n8080_o;
  wire n8082_o;
  wire n8083_o;
  wire [7:0] n8085_o;
  wire n8087_o;
  wire n8088_o;
  wire n8091_o;
  wire n8093_o;
  wire n8099_o;
  wire n8102_o;
  wire n8104_o;
  wire n8106_o;
  wire n8108_o;
  wire n8110_o;
  wire n8112_o;
  wire n8114_o;
  wire n8116_o;
  wire n8118_o;
  wire n8120_o;
  wire n8122_o;
  wire [10:0] n8123_o;
  reg [7:0] n8129_o;
  wire n8131_o;
  wire [15:0] n8134_o;
  wire n8136_o;
  wire n8138_o;
  wire n8140_o;
  wire [3:0] n8141_o;
  reg [15:0] n8142_o;
  wire n8144_o;
  wire n8145_o;
  wire n8147_o;
  wire [1:0] n8148_o;
  reg n8149_o;
  wire n8215_o;
  wire [16:0] n8216_o;
  wire [16:0] n8217_o;
  wire [16:0] n8218_o;
  wire [15:0] n8219_o;
  wire n8221_o;
  localparam [7:0] n8222_o = 8'b00000000;
  wire n8224_o;
  wire [4:0] n8225_o;
  wire [2:0] n8226_o;
  wire n8228_o;
  wire [15:0] n8229_o;
  wire [15:0] n8230_o;
  wire [15:0] n8231_o;
  wire n8233_o;
  wire n8235_o;
  wire n8237_o;
  wire n8239_o;
  wire [15:0] n8240_o;
  wire [15:0] n8241_o;
  wire n8243_o;
  wire [8:0] n8244_o;
  wire [7:0] n8245_o;
  wire [7:0] n8246_o;
  wire [7:0] n8247_o;
  wire [7:0] n8248_o;
  wire [7:0] n8249_o;
  wire [7:0] n8250_o;
  reg [7:0] n8251_o;
  wire [2:0] n8252_o;
  wire [2:0] n8253_o;
  wire [2:0] n8254_o;
  wire [2:0] n8255_o;
  wire [2:0] n8256_o;
  wire [2:0] n8257_o;
  wire [2:0] n8258_o;
  wire [2:0] n8259_o;
  wire [2:0] n8260_o;
  reg [2:0] n8261_o;
  wire [4:0] n8262_o;
  wire [4:0] n8263_o;
  wire [4:0] n8264_o;
  wire [4:0] n8265_o;
  wire [4:0] n8266_o;
  wire [4:0] n8267_o;
  wire [4:0] n8268_o;
  wire [4:0] n8269_o;
  wire [4:0] n8270_o;
  reg [4:0] n8271_o;
  wire n8293_o;
  wire n8294_o;
  wire n8295_o;
  wire n8296_o;
  wire n8297_o;
  wire n8298_o;
  wire n8299_o;
  wire n8300_o;
  wire n8301_o;
  wire n8302_o;
  wire n8303_o;
  wire n8304_o;
  wire n8305_o;
  wire n8306_o;
  wire n8307_o;
  wire n8308_o;
  wire n8309_o;
  wire n8310_o;
  wire n8311_o;
  wire n8312_o;
  wire n8313_o;
  wire n8314_o;
  wire n8315_o;
  wire n8316_o;
  wire n8317_o;
  wire n8318_o;
  wire n8319_o;
  wire n8320_o;
  wire n8321_o;
  wire n8322_o;
  wire n8323_o;
  wire n8324_o;
  wire n8325_o;
  wire n8326_o;
  wire n8328_o;
  wire n8329_o;
  wire n8330_o;
  wire [7:0] n8333_o;
  wire [7:0] n8336_o;
  wire n8338_o;
  wire n8340_o;
  wire n8341_o;
  wire [7:0] n8344_o;
  reg [7:0] n8345_o;
  wire [7:0] n8346_o;
  wire n8348_o;
  wire n8350_o;
  wire n8351_o;
  wire n8352_o;
  wire n8354_o;
  wire [31:0] n8355_o;
  wire n8357_o;
  wire [7:0] n8358_o;
  wire n8360_o;
  wire n8361_o;
  wire n8362_o;
  wire n8364_o;
  wire n8365_o;
  wire n8366_o;
  wire [7:0] n8369_o;
  wire n8371_o;
  wire [31:0] n8372_o;
  wire n8374_o;
  wire [7:0] n8377_o;
  wire [7:0] n8378_o;
  wire [7:0] n8381_o;
  wire [7:0] n8382_o;
  wire [7:0] n8383_o;
  wire n8385_o;
  wire [1:0] n8386_o;
  reg [7:0] n8387_o;
  wire n8388_o;
  wire [31:0] n8389_o;
  wire n8391_o;
  wire n8393_o;
  wire n8395_o;
  wire [3:0] n8396_o;
  wire n8397_o;
  wire n8399_o;
  wire n8401_o;
  wire n8403_o;
  wire n8405_o;
  wire n8407_o;
  wire n8409_o;
  wire n8411_o;
  wire n8413_o;
  wire n8415_o;
  wire n8417_o;
  wire n8419_o;
  wire n8421_o;
  wire n8423_o;
  wire n8425_o;
  wire n8427_o;
  wire n8429_o;
  wire [6:0] n8430_o;
  wire n8432_o;
  wire n8434_o;
  wire n8436_o;
  wire [21:0] n8437_o;
  reg n8440_o;
  reg n8446_o;
  reg n8447_o;
  reg [7:0] n8448_o;
  reg [1:0] n8453_o;
  reg [7:0] n8454_o;
  reg [7:0] n8455_o;
  reg [7:0] n8456_o;
  reg [3:0] n8457_o;
  wire n8458_o;
  wire n8459_o;
  wire n8460_o;
  wire n8461_o;
  wire [7:0] n8462_o;
  reg [7:0] n8463_o;
  reg [7:0] n8464_o;
  reg [7:0] n8465_o;
  wire [5:0] n8466_o;
  wire [7:0] n8467_o;
  reg [7:0] n8468_o;
  reg [7:0] n8469_o;
  reg [7:0] n8470_o;
  reg [7:0] n8471_o;
  reg [7:0] n8472_o;
  reg [7:0] n8473_o;
  wire [6:0] n8474_o;
  reg [6:0] n8475_o;
  reg [7:0] n8476_o;
  reg [7:0] n8477_o;
  reg [7:0] n8478_o;
  reg [7:0] n8479_o;
  wire [3:0] n8480_o;
  wire n8482_o;
  wire [3:0] n8483_o;
  wire n8488_o;
  wire n8490_o;
  wire n8492_o;
  wire n8494_o;
  wire n8496_o;
  wire n8498_o;
  wire n8500_o;
  wire n8502_o;
  wire [7:0] n8503_o;
  wire [7:0] n8504_o;
  wire [7:0] n8505_o;
  wire [7:0] n8506_o;
  wire [7:0] n8507_o;
  wire [7:0] n8508_o;
  wire [7:0] n8509_o;
  wire [7:0] n8510_o;
  wire [7:0] n8511_o;
  wire [7:0] n8512_o;
  wire [7:0] n8513_o;
  wire [7:0] n8514_o;
  wire [7:0] n8515_o;
  wire [7:0] n8516_o;
  wire [7:0] n8517_o;
  wire [7:0] n8518_o;
  wire [7:0] n8519_o;
  wire [7:0] n8520_o;
  wire [7:0] n8521_o;
  wire [7:0] n8522_o;
  wire [7:0] n8523_o;
  wire [7:0] n8524_o;
  wire [7:0] n8525_o;
  wire [7:0] n8526_o;
  wire [7:0] n8527_o;
  wire [7:0] n8528_o;
  wire [7:0] n8529_o;
  wire [7:0] n8530_o;
  wire [7:0] n8531_o;
  wire [7:0] n8532_o;
  wire [7:0] n8533_o;
  wire [7:0] n8534_o;
  wire [7:0] n8535_o;
  wire [7:0] n8536_o;
  wire [7:0] n8537_o;
  wire [7:0] n8538_o;
  wire [127:0] n8539_o;
  wire [7:0] n8540_o;
  wire [7:0] n8541_o;
  wire [7:0] n8542_o;
  wire [7:0] n8543_o;
  wire [7:0] n8544_o;
  wire [7:0] n8545_o;
  wire [7:0] n8546_o;
  wire [7:0] n8547_o;
  wire n8549_o;
  wire n8551_o;
  wire [127:0] n8552_o;
  wire [7:0] n8553_o;
  wire [7:0] n8554_o;
  wire [7:0] n8555_o;
  wire [7:0] n8556_o;
  wire [7:0] n8557_o;
  wire [7:0] n8558_o;
  wire [7:0] n8559_o;
  wire [7:0] n8560_o;
  wire n8561_o;
  wire [7:0] n8562_o;
  wire [1:0] n8563_o;
  wire [7:0] n8564_o;
  wire [7:0] n8565_o;
  wire [7:0] n8566_o;
  wire [3:0] n8567_o;
  wire n8568_o;
  wire n8569_o;
  wire n8570_o;
  wire n8571_o;
  wire [7:0] n8572_o;
  wire [7:0] n8573_o;
  wire [7:0] n8574_o;
  wire [7:0] n8575_o;
  wire [5:0] n8576_o;
  wire [7:0] n8577_o;
  wire [7:0] n8578_o;
  wire [7:0] n8579_o;
  wire [7:0] n8580_o;
  wire [7:0] n8581_o;
  wire [7:0] n8582_o;
  wire [7:0] n8583_o;
  wire [6:0] n8584_o;
  wire [6:0] n8585_o;
  wire [7:0] n8586_o;
  wire [7:0] n8587_o;
  wire [7:0] n8588_o;
  wire [7:0] n8589_o;
  wire n8591_o;
  wire n8593_o;
  wire n8594_o;
  wire n8595_o;
  wire n8596_o;
  wire n8598_o;
  wire n8599_o;
  wire n8600_o;
  wire n8602_o;
  wire n8604_o;
  wire n8605_o;
  wire n8607_o;
  wire n8608_o;
  wire n8610_o;
  wire n8611_o;
  wire n8613_o;
  wire n8614_o;
  wire n8615_o;
  wire n8616_o;
  wire [3:0] n8617_o;
  wire [2:0] n8618_o;
  wire n8623_o;
  wire [2:0] n8624_o;
  wire n8627_o;
  wire n8628_o;
  wire n8629_o;
  wire n8630_o;
  wire [7:0] n8631_o;
  wire n8634_o;
  wire [2:0] n8635_o;
  wire n8640_o;
  wire [2:0] n8641_o;
  wire [5:0] n8644_o;
  wire [7:0] n8645_o;
  wire n8648_o;
  wire [2:0] n8649_o;
  wire n8654_o;
  wire [2:0] n8655_o;
  wire n8660_o;
  wire [2:0] n8661_o;
  wire n8666_o;
  wire [2:0] n8667_o;
  wire n8672_o;
  wire [2:0] n8673_o;
  wire n8675_o;
  wire n8677_o;
  wire n8679_o;
  wire n8681_o;
  wire n8683_o;
  wire n8685_o;
  wire n8687_o;
  wire n8689_o;
  wire [7:0] n8690_o;
  wire n8691_o;
  reg n8692_o;
  wire n8693_o;
  reg n8694_o;
  wire n8695_o;
  reg n8696_o;
  wire n8697_o;
  reg n8698_o;
  wire n8699_o;
  reg n8700_o;
  wire n8701_o;
  reg n8702_o;
  wire n8703_o;
  reg n8704_o;
  wire n8706_o;
  wire [2:0] n8707_o;
  wire n8712_o;
  wire [2:0] n8713_o;
  wire n8718_o;
  wire [10:0] n8719_o;
  reg [7:0] n8720_o;
  wire n8721_o;
  wire n8722_o;
  wire n8723_o;
  wire n8724_o;
  wire [7:0] n8725_o;
  reg [7:0] n8726_o;
  reg [7:0] n8727_o;
  wire [5:0] n8728_o;
  wire [7:0] n8729_o;
  reg [7:0] n8730_o;
  reg [7:0] n8731_o;
  reg [7:0] n8732_o;
  reg [7:0] n8733_o;
  reg [7:0] n8734_o;
  wire n8735_o;
  reg n8736_o;
  wire n8737_o;
  reg n8738_o;
  wire n8739_o;
  reg n8740_o;
  wire n8741_o;
  reg n8742_o;
  wire n8743_o;
  reg n8744_o;
  wire n8745_o;
  reg n8746_o;
  wire n8747_o;
  reg n8748_o;
  reg [7:0] n8749_o;
  reg [7:0] n8750_o;
  wire [3:0] n8751_o;
  wire [2:0] n8754_o;
  wire [127:0] n8759_o;
  wire [7:0] n8760_o;
  wire n8761_o;
  wire n8762_o;
  wire n8763_o;
  wire n8764_o;
  wire [7:0] n8765_o;
  wire [7:0] n8766_o;
  wire [7:0] n8767_o;
  wire [5:0] n8768_o;
  wire [7:0] n8769_o;
  wire [7:0] n8770_o;
  wire [7:0] n8771_o;
  wire [7:0] n8772_o;
  wire [7:0] n8773_o;
  wire [7:0] n8774_o;
  wire [6:0] n8775_o;
  wire [6:0] n8776_o;
  wire [6:0] n8777_o;
  wire [7:0] n8778_o;
  wire [7:0] n8779_o;
  wire [127:0] n8780_o;
  wire n8781_o;
  wire n8782_o;
  wire n8783_o;
  wire n8784_o;
  wire n8785_o;
  wire [7:0] n8786_o;
  wire [7:0] n8787_o;
  wire n8788_o;
  wire [5:0] n8789_o;
  wire [7:0] n8790_o;
  wire [7:0] n8791_o;
  wire n8792_o;
  wire n8793_o;
  wire n8794_o;
  wire n8795_o;
  wire [5:0] n8796_o;
  wire [5:0] n8797_o;
  wire [5:0] n8798_o;
  wire n8799_o;
  wire n8800_o;
  wire n8801_o;
  wire n8802_o;
  wire n8804_o;
  wire n8805_o;
  wire n8807_o;
  wire n8809_o;
  wire n8810_o;
  wire n8812_o;
  wire n8813_o;
  wire n8816_o;
  wire n8818_o;
  wire n8819_o;
  wire [1:0] n8820_o;
  wire n8821_o;
  reg n8822_o;
  wire n8823_o;
  reg n8824_o;
  reg [7:0] n8825_o;
  reg [7:0] n8826_o;
  wire n8828_o;
  wire [5:0] n8829_o;
  reg n8831_o;
  reg n8834_o;
  reg [127:0] n8836_o;
  reg [7:0] n8837_o;
  reg [7:0] n8838_o;
  reg [7:0] n8839_o;
  reg [7:0] n8840_o;
  reg [7:0] n8841_o;
  reg [7:0] n8842_o;
  reg [7:0] n8843_o;
  reg [7:0] n8844_o;
  reg n8845_o;
  reg [7:0] n8846_o;
  reg [1:0] n8847_o;
  reg [7:0] n8848_o;
  reg [7:0] n8849_o;
  reg [7:0] n8850_o;
  reg [7:0] n8851_o;
  reg [3:0] n8852_o;
  wire n8853_o;
  wire n8854_o;
  wire n8855_o;
  wire n8856_o;
  wire [7:0] n8857_o;
  reg [7:0] n8858_o;
  reg [7:0] n8859_o;
  reg [7:0] n8860_o;
  wire [5:0] n8861_o;
  wire [7:0] n8862_o;
  reg [7:0] n8863_o;
  reg [7:0] n8864_o;
  reg [7:0] n8865_o;
  reg [7:0] n8866_o;
  reg [7:0] n8867_o;
  reg [7:0] n8868_o;
  wire n8869_o;
  wire n8870_o;
  wire n8871_o;
  reg n8872_o;
  wire n8873_o;
  wire n8874_o;
  wire n8875_o;
  reg n8876_o;
  wire [2:0] n8877_o;
  wire [2:0] n8878_o;
  wire [2:0] n8879_o;
  reg [2:0] n8880_o;
  wire n8881_o;
  wire n8882_o;
  wire n8883_o;
  reg n8884_o;
  wire n8885_o;
  wire n8886_o;
  reg n8887_o;
  reg [7:0] n8888_o;
  reg [7:0] n8889_o;
  reg [7:0] n8890_o;
  reg [7:0] n8891_o;
  wire [7:0] n8920_o;
  wire n8928_o;
  wire [127:0] n8933_o;
  wire [7:0] n8996_o;
  reg [7:0] n8997_q;
  wire [15:0] n8998_o;
  reg [15:0] n8999_q;
  wire n9000_o;
  reg n9001_q;
  wire n9002_o;
  wire [7:0] n9003_o;
  reg [7:0] n9004_q;
  wire [127:0] n9005_o;
  reg [127:0] n9006_q;
  wire [7:0] n9007_o;
  reg [7:0] n9008_q;
  wire [7:0] n9009_o;
  reg [7:0] n9010_q;
  wire [7:0] n9011_o;
  reg [7:0] n9012_q;
  wire [7:0] n9013_o;
  reg [7:0] n9014_q;
  wire [7:0] n9015_o;
  reg [7:0] n9016_q;
  wire [7:0] n9017_o;
  reg [7:0] n9018_q;
  wire [7:0] n9019_o;
  reg [7:0] n9020_q;
  wire [7:0] n9021_o;
  reg [7:0] n9022_q;
  wire [2:0] n9023_o;
  reg [2:0] n9024_q;
  wire n9025_o;
  wire n9026_o;
  reg n9027_q;
  wire n9028_o;
  wire n9029_o;
  reg n9030_q;
  wire n9031_o;
  wire n9032_o;
  reg n9033_q;
  wire n9034_o;
  wire n9035_o;
  reg n9036_q;
  wire n9037_o;
  wire n9038_o;
  reg n9039_q;
  wire n9040_o;
  wire n9041_o;
  reg n9042_q;
  wire n9043_o;
  wire n9044_o;
  reg n9045_q;
  wire n9046_o;
  reg n9047_q;
  wire n9048_o;
  reg n9049_q;
  wire [7:0] n9050_o;
  reg [7:0] n9051_q;
  wire [1:0] n9052_o;
  reg [1:0] n9053_q;
  wire n9054_o;
  reg n9055_q;
  wire n9056_o;
  reg n9057_q;
  wire n9058_o;
  reg n9059_q;
  wire n9060_o;
  reg n9061_q;
  wire n9062_o;
  reg n9063_q;
  wire n9064_o;
  reg n9065_q;
  wire n9066_o;
  reg n9067_q;
  wire n9068_o;
  reg n9069_q;
  wire n9070_o;
  reg n9071_q;
  wire n9072_o;
  reg n9073_q;
  wire n9074_o;
  reg n9075_q;
  wire n9076_o;
  reg n9077_q;
  wire n9078_o;
  reg n9079_q;
  wire n9080_o;
  reg n9081_q;
  wire [7:0] n9084_o;
  reg [7:0] n9085_q;
  wire [7:0] n9086_o;
  reg [7:0] n9087_q;
  wire [7:0] n9088_o;
  reg [7:0] n9089_q;
  wire [7:0] n9090_o;
  reg [7:0] n9091_q;
  wire [15:0] n9092_o;
  reg [15:0] n9093_q;
  wire [15:0] n9094_o;
  wire [7:0] n9095_o;
  wire [7:0] n9096_o;
  reg [7:0] n9097_q;
  wire [7:0] n9098_o;
  reg [7:0] n9099_q;
  wire [7:0] n9100_o;
  reg [7:0] n9101_q;
  wire [7:0] n9102_o;
  reg [7:0] n9103_q;
  wire [7:0] n9104_o;
  reg [7:0] n9105_q;
  wire [3:0] n9106_o;
  reg [3:0] n9107_q;
  wire [7:0] n9108_o;
  reg [7:0] n9109_q;
  wire [7:0] n9110_o;
  reg [7:0] n9111_q;
  wire [7:0] n9112_o;
  reg [7:0] n9113_q;
  wire [7:0] n9114_o;
  reg [7:0] n9115_q;
  wire [7:0] n9116_o;
  reg [7:0] n9117_q;
  wire [7:0] n9118_o;
  reg [7:0] n9119_q;
  wire [7:0] n9120_o;
  reg [7:0] n9121_q;
  wire [7:0] n9122_o;
  reg [7:0] n9123_q;
  wire [7:0] n9124_o;
  reg [7:0] n9125_q;
  wire [7:0] n9126_o;
  reg [7:0] n9127_q;
  wire [7:0] n9128_o;
  reg [7:0] n9129_q;
  wire [7:0] n9130_o;
  reg [7:0] n9131_q;
  wire [7:0] n9132_o;
  reg [7:0] n9133_q;
  wire [7:0] n9134_o;
  reg [7:0] n9135_q;
  wire [1:0] n9136_o;
  wire n9137_o;
  reg n9138_q;
  wire [5:0] n9139_o;
  wire n9140_o;
  reg n9141_q;
  wire [15:0] n9142_o;
  wire [7:0] n9144_o;
  wire [7:0] n9145_o;
  wire [7:0] n9146_o;
  wire [7:0] n9147_o;
  wire [7:0] n9148_o;
  wire [7:0] n9149_o;
  wire [7:0] n9150_o;
  wire [7:0] n9151_o;
  wire [7:0] n9152_o;
  wire [7:0] n9153_o;
  wire [7:0] n9154_o;
  wire [7:0] n9155_o;
  wire [7:0] n9156_o;
  wire [7:0] n9157_o;
  wire [7:0] n9158_o;
  wire [7:0] n9159_o;
  wire [1:0] n9160_o;
  reg [7:0] n9161_o;
  wire [1:0] n9162_o;
  reg [7:0] n9163_o;
  wire [1:0] n9164_o;
  reg [7:0] n9165_o;
  wire [1:0] n9166_o;
  reg [7:0] n9167_o;
  wire [1:0] n9168_o;
  reg [7:0] n9169_o;
  wire n9170_o;
  wire n9171_o;
  wire n9172_o;
  wire n9173_o;
  wire n9174_o;
  wire n9175_o;
  wire n9176_o;
  wire n9177_o;
  wire [1:0] n9178_o;
  reg n9179_o;
  wire [1:0] n9180_o;
  reg n9181_o;
  wire n9182_o;
  wire n9183_o;
  wire n9184_o;
  wire n9185_o;
  wire n9186_o;
  wire n9187_o;
  wire n9188_o;
  wire n9189_o;
  wire n9190_o;
  wire n9191_o;
  wire [1:0] n9192_o;
  reg n9193_o;
  wire [1:0] n9194_o;
  reg n9195_o;
  wire n9196_o;
  wire n9197_o;
  wire n9198_o;
  wire n9199_o;
  wire n9200_o;
  wire n9201_o;
  wire n9202_o;
  wire n9203_o;
  wire n9204_o;
  wire n9205_o;
  wire [1:0] n9206_o;
  reg n9207_o;
  wire [1:0] n9208_o;
  reg n9209_o;
  wire n9210_o;
  wire n9211_o;
  wire n9212_o;
  wire n9213_o;
  wire n9214_o;
  wire n9215_o;
  wire n9216_o;
  wire n9217_o;
  wire n9218_o;
  wire n9219_o;
  wire [1:0] n9220_o;
  reg n9221_o;
  wire [1:0] n9222_o;
  reg n9223_o;
  wire n9224_o;
  wire n9225_o;
  wire n9226_o;
  wire n9227_o;
  wire n9228_o;
  wire n9229_o;
  wire n9230_o;
  wire n9231_o;
  wire n9232_o;
  wire n9233_o;
  wire [1:0] n9234_o;
  reg n9235_o;
  wire [1:0] n9236_o;
  reg n9237_o;
  wire n9238_o;
  wire n9239_o;
  wire n9240_o;
  wire n9241_o;
  wire n9242_o;
  wire n9243_o;
  wire n9244_o;
  wire n9245_o;
  wire n9246_o;
  wire n9247_o;
  wire [1:0] n9248_o;
  reg n9249_o;
  wire [1:0] n9250_o;
  reg n9251_o;
  wire n9252_o;
  wire n9253_o;
  wire n9254_o;
  wire n9255_o;
  wire n9256_o;
  wire n9257_o;
  wire n9258_o;
  wire n9259_o;
  wire n9260_o;
  wire n9261_o;
  wire [1:0] n9262_o;
  reg n9263_o;
  wire [1:0] n9264_o;
  reg n9265_o;
  wire n9266_o;
  wire n9267_o;
  wire n9268_o;
  wire n9269_o;
  wire n9270_o;
  wire n9271_o;
  wire n9272_o;
  wire n9273_o;
  wire n9274_o;
  wire n9275_o;
  wire [1:0] n9276_o;
  reg n9277_o;
  wire [1:0] n9278_o;
  reg n9279_o;
  wire n9280_o;
  wire n9281_o;
  wire n9282_o;
  wire n9283_o;
  wire n9284_o;
  wire n9285_o;
  wire n9286_o;
  wire n9287_o;
  wire n9288_o;
  wire n9289_o;
  wire [1:0] n9290_o;
  reg n9291_o;
  wire [1:0] n9292_o;
  reg n9293_o;
  wire n9294_o;
  wire n9295_o;
  wire n9296_o;
  wire n9297_o;
  wire n9298_o;
  wire n9299_o;
  wire n9300_o;
  wire n9301_o;
  wire n9302_o;
  wire n9303_o;
  wire [1:0] n9304_o;
  reg n9305_o;
  wire [1:0] n9306_o;
  reg n9307_o;
  wire n9308_o;
  wire n9309_o;
  wire n9310_o;
  wire n9311_o;
  wire n9312_o;
  wire n9313_o;
  wire n9314_o;
  wire n9315_o;
  wire n9316_o;
  wire n9317_o;
  wire [1:0] n9318_o;
  reg n9319_o;
  wire [1:0] n9320_o;
  reg n9321_o;
  wire n9322_o;
  wire n9323_o;
  wire n9324_o;
  wire n9325_o;
  wire n9326_o;
  wire n9327_o;
  wire n9328_o;
  wire n9329_o;
  wire n9330_o;
  wire n9331_o;
  wire n9332_o;
  wire n9333_o;
  wire n9334_o;
  wire n9335_o;
  wire n9336_o;
  wire n9337_o;
  wire n9338_o;
  wire n9339_o;
  wire n9340_o;
  wire n9341_o;
  wire n9342_o;
  wire n9343_o;
  wire n9344_o;
  wire n9345_o;
  wire n9346_o;
  wire n9347_o;
  wire n9348_o;
  wire n9349_o;
  wire n9350_o;
  wire n9351_o;
  wire n9352_o;
  wire n9353_o;
  wire n9354_o;
  wire n9355_o;
  wire n9356_o;
  wire n9357_o;
  wire n9358_o;
  wire n9359_o;
  wire n9360_o;
  wire n9361_o;
  wire n9362_o;
  wire n9363_o;
  wire n9364_o;
  wire n9365_o;
  wire n9366_o;
  wire n9367_o;
  wire n9368_o;
  wire n9369_o;
  wire n9370_o;
  wire n9371_o;
  wire n9372_o;
  wire n9373_o;
  wire n9374_o;
  wire n9375_o;
  wire n9376_o;
  wire n9377_o;
  wire n9378_o;
  wire n9379_o;
  wire n9380_o;
  wire n9381_o;
  wire n9382_o;
  wire n9383_o;
  wire n9384_o;
  wire n9385_o;
  wire n9386_o;
  wire n9387_o;
  wire n9388_o;
  wire n9389_o;
  wire n9390_o;
  wire n9391_o;
  wire n9392_o;
  wire n9393_o;
  wire n9394_o;
  wire n9395_o;
  wire n9396_o;
  wire n9397_o;
  wire n9398_o;
  wire n9399_o;
  wire n9400_o;
  wire n9401_o;
  wire n9402_o;
  wire n9403_o;
  wire n9404_o;
  wire n9405_o;
  wire n9406_o;
  wire n9407_o;
  wire n9408_o;
  wire n9409_o;
  wire n9410_o;
  wire n9411_o;
  wire n9412_o;
  wire n9413_o;
  wire n9414_o;
  wire n9415_o;
  wire n9416_o;
  wire n9417_o;
  wire n9418_o;
  wire n9419_o;
  wire n9420_o;
  wire n9421_o;
  wire n9422_o;
  wire n9423_o;
  wire n9424_o;
  wire n9425_o;
  wire n9426_o;
  wire n9427_o;
  wire n9428_o;
  wire n9429_o;
  wire n9430_o;
  wire n9431_o;
  wire n9432_o;
  wire n9433_o;
  wire n9434_o;
  wire n9435_o;
  wire n9436_o;
  wire n9437_o;
  wire n9438_o;
  wire n9439_o;
  wire n9440_o;
  wire n9441_o;
  wire n9442_o;
  wire n9443_o;
  wire n9444_o;
  wire n9445_o;
  wire n9446_o;
  wire n9447_o;
  wire n9448_o;
  wire n9449_o;
  wire n9450_o;
  wire n9451_o;
  wire [6:0] n9452_o;
  wire [1:0] n9453_o;
  reg n9454_o;
  wire [1:0] n9455_o;
  reg n9456_o;
  wire [1:0] n9457_o;
  reg n9458_o;
  wire [1:0] n9459_o;
  reg n9460_o;
  wire [1:0] n9461_o;
  reg n9462_o;
  wire [1:0] n9463_o;
  reg n9464_o;
  wire [1:0] n9465_o;
  reg n9466_o;
  wire [1:0] n9467_o;
  reg n9468_o;
  wire [1:0] n9469_o;
  reg n9470_o;
  wire [1:0] n9471_o;
  reg n9472_o;
  wire [1:0] n9473_o;
  reg n9474_o;
  wire [1:0] n9475_o;
  reg n9476_o;
  wire [1:0] n9477_o;
  reg n9478_o;
  wire [1:0] n9479_o;
  reg n9480_o;
  wire [1:0] n9481_o;
  reg n9482_o;
  wire [1:0] n9483_o;
  reg n9484_o;
  wire [1:0] n9485_o;
  reg n9486_o;
  wire [1:0] n9487_o;
  reg n9488_o;
  wire [1:0] n9489_o;
  reg n9490_o;
  wire [1:0] n9491_o;
  reg n9492_o;
  wire [1:0] n9493_o;
  reg n9494_o;
  wire [1:0] n9495_o;
  reg n9496_o;
  wire [1:0] n9497_o;
  reg n9498_o;
  wire [1:0] n9499_o;
  reg n9500_o;
  wire [1:0] n9501_o;
  reg n9502_o;
  wire [1:0] n9503_o;
  reg n9504_o;
  wire [1:0] n9505_o;
  reg n9506_o;
  wire [1:0] n9507_o;
  reg n9508_o;
  wire [1:0] n9509_o;
  reg n9510_o;
  wire [1:0] n9511_o;
  reg n9512_o;
  wire [1:0] n9513_o;
  reg n9514_o;
  wire [1:0] n9515_o;
  reg n9516_o;
  wire [1:0] n9517_o;
  reg n9518_o;
  wire [1:0] n9519_o;
  reg n9520_o;
  wire [1:0] n9521_o;
  reg n9522_o;
  wire [1:0] n9523_o;
  reg n9524_o;
  wire [1:0] n9525_o;
  reg n9526_o;
  wire [1:0] n9527_o;
  reg n9528_o;
  wire [1:0] n9529_o;
  reg n9530_o;
  wire [1:0] n9531_o;
  reg n9532_o;
  wire [1:0] n9533_o;
  reg n9534_o;
  wire [1:0] n9535_o;
  reg n9536_o;
  wire n9537_o;
  wire n9538_o;
  wire n9539_o;
  wire n9540_o;
  wire n9541_o;
  wire n9542_o;
  wire n9543_o;
  wire n9544_o;
  wire n9545_o;
  wire n9546_o;
  wire n9547_o;
  wire n9548_o;
  wire n9549_o;
  wire n9550_o;
  wire n9551_o;
  wire n9552_o;
  wire n9553_o;
  wire n9554_o;
  wire n9555_o;
  wire n9556_o;
  wire n9557_o;
  wire n9558_o;
  wire n9559_o;
  wire n9560_o;
  wire n9561_o;
  wire n9562_o;
  wire n9563_o;
  wire n9564_o;
  wire n9565_o;
  wire n9566_o;
  wire n9567_o;
  wire n9568_o;
  wire n9569_o;
  wire n9570_o;
  wire n9571_o;
  wire n9572_o;
  wire n9573_o;
  wire n9574_o;
  wire [7:0] n9575_o;
  wire [7:0] n9576_o;
  wire [7:0] n9577_o;
  wire [7:0] n9578_o;
  wire [7:0] n9579_o;
  wire [7:0] n9580_o;
  wire [7:0] n9581_o;
  wire [7:0] n9582_o;
  wire [7:0] n9583_o;
  wire [7:0] n9584_o;
  wire [7:0] n9585_o;
  wire [7:0] n9586_o;
  wire [7:0] n9587_o;
  wire [7:0] n9588_o;
  wire [7:0] n9589_o;
  wire [7:0] n9590_o;
  wire [7:0] n9591_o;
  wire [7:0] n9592_o;
  wire [7:0] n9593_o;
  wire [7:0] n9594_o;
  wire [7:0] n9595_o;
  wire [7:0] n9596_o;
  wire [7:0] n9597_o;
  wire [7:0] n9598_o;
  wire [7:0] n9599_o;
  wire [7:0] n9600_o;
  wire [7:0] n9601_o;
  wire [7:0] n9602_o;
  wire [7:0] n9603_o;
  wire [7:0] n9604_o;
  wire [7:0] n9605_o;
  wire [7:0] n9606_o;
  wire [127:0] n9607_o;
  wire n9608_o;
  wire n9609_o;
  wire n9610_o;
  wire n9611_o;
  wire n9612_o;
  wire n9613_o;
  wire n9614_o;
  wire n9615_o;
  wire n9616_o;
  wire n9617_o;
  wire n9618_o;
  wire n9619_o;
  wire n9620_o;
  wire n9621_o;
  wire n9622_o;
  wire n9623_o;
  wire n9624_o;
  wire n9625_o;
  wire n9626_o;
  wire n9627_o;
  wire n9628_o;
  wire n9629_o;
  wire n9630_o;
  wire n9631_o;
  wire n9632_o;
  wire n9633_o;
  wire n9634_o;
  wire n9635_o;
  wire n9636_o;
  wire n9637_o;
  wire n9638_o;
  wire n9639_o;
  wire n9640_o;
  wire n9641_o;
  wire [7:0] n9642_o;
  wire n9643_o;
  wire n9644_o;
  wire n9645_o;
  wire n9646_o;
  wire n9647_o;
  wire n9648_o;
  wire n9649_o;
  wire n9650_o;
  wire n9651_o;
  wire n9652_o;
  wire n9653_o;
  wire n9654_o;
  wire n9655_o;
  wire n9656_o;
  wire n9657_o;
  wire n9658_o;
  wire n9659_o;
  wire n9660_o;
  wire n9661_o;
  wire n9662_o;
  wire n9663_o;
  wire n9664_o;
  wire n9665_o;
  wire n9666_o;
  wire n9667_o;
  wire n9668_o;
  wire n9669_o;
  wire n9670_o;
  wire n9671_o;
  wire n9672_o;
  wire n9673_o;
  wire n9674_o;
  wire n9675_o;
  wire n9676_o;
  wire [7:0] n9677_o;
  wire n9678_o;
  wire n9679_o;
  wire n9680_o;
  wire n9681_o;
  wire n9682_o;
  wire n9683_o;
  wire n9684_o;
  wire n9685_o;
  wire n9686_o;
  wire n9687_o;
  wire n9688_o;
  wire n9689_o;
  wire n9690_o;
  wire n9691_o;
  wire n9692_o;
  wire n9693_o;
  wire n9694_o;
  wire n9695_o;
  wire n9696_o;
  wire n9697_o;
  wire n9698_o;
  wire n9699_o;
  wire n9700_o;
  wire n9701_o;
  wire n9702_o;
  wire n9703_o;
  wire n9704_o;
  wire n9705_o;
  wire n9706_o;
  wire n9707_o;
  wire n9708_o;
  wire n9709_o;
  wire n9710_o;
  wire n9711_o;
  wire [7:0] n9712_o;
  wire n9713_o;
  wire n9714_o;
  wire n9715_o;
  wire n9716_o;
  wire n9717_o;
  wire n9718_o;
  wire n9719_o;
  wire n9720_o;
  wire n9721_o;
  wire n9722_o;
  wire n9723_o;
  wire n9724_o;
  wire n9725_o;
  wire n9726_o;
  wire n9727_o;
  wire n9728_o;
  wire n9729_o;
  wire n9730_o;
  wire n9731_o;
  wire n9732_o;
  wire n9733_o;
  wire n9734_o;
  wire n9735_o;
  wire n9736_o;
  wire n9737_o;
  wire n9738_o;
  wire n9739_o;
  wire n9740_o;
  wire n9741_o;
  wire n9742_o;
  wire n9743_o;
  wire n9744_o;
  wire n9745_o;
  wire n9746_o;
  wire [7:0] n9747_o;
  wire n9748_o;
  wire n9749_o;
  wire n9750_o;
  wire n9751_o;
  wire n9752_o;
  wire n9753_o;
  wire n9754_o;
  wire n9755_o;
  wire n9756_o;
  wire n9757_o;
  wire n9758_o;
  wire n9759_o;
  wire n9760_o;
  wire n9761_o;
  wire n9762_o;
  wire n9763_o;
  wire n9764_o;
  wire n9765_o;
  wire n9766_o;
  wire n9767_o;
  wire n9768_o;
  wire n9769_o;
  wire n9770_o;
  wire n9771_o;
  wire n9772_o;
  wire n9773_o;
  wire n9774_o;
  wire n9775_o;
  wire n9776_o;
  wire n9777_o;
  wire n9778_o;
  wire n9779_o;
  wire n9780_o;
  wire n9781_o;
  wire [7:0] n9782_o;
  wire n9783_o;
  wire n9784_o;
  wire n9785_o;
  wire n9786_o;
  wire n9787_o;
  wire n9788_o;
  wire n9789_o;
  wire n9790_o;
  wire n9791_o;
  wire n9792_o;
  wire n9793_o;
  wire n9794_o;
  wire n9795_o;
  wire n9796_o;
  wire n9797_o;
  wire n9798_o;
  wire n9799_o;
  wire n9800_o;
  wire n9801_o;
  wire n9802_o;
  wire n9803_o;
  wire n9804_o;
  wire n9805_o;
  wire n9806_o;
  wire n9807_o;
  wire n9808_o;
  wire n9809_o;
  wire n9810_o;
  wire n9811_o;
  wire n9812_o;
  wire n9813_o;
  wire n9814_o;
  wire n9815_o;
  wire n9816_o;
  wire [7:0] n9817_o;
  wire n9818_o;
  wire n9819_o;
  wire n9820_o;
  wire n9821_o;
  wire n9822_o;
  wire n9823_o;
  wire n9824_o;
  wire n9825_o;
  wire n9826_o;
  wire n9827_o;
  wire n9828_o;
  wire n9829_o;
  wire n9830_o;
  wire n9831_o;
  wire n9832_o;
  wire n9833_o;
  wire n9834_o;
  wire n9835_o;
  wire n9836_o;
  wire n9837_o;
  wire n9838_o;
  wire n9839_o;
  wire n9840_o;
  wire n9841_o;
  wire n9842_o;
  wire n9843_o;
  wire n9844_o;
  wire n9845_o;
  wire n9846_o;
  wire n9847_o;
  wire n9848_o;
  wire n9849_o;
  wire n9850_o;
  wire n9851_o;
  wire [7:0] n9852_o;
  wire n9853_o;
  wire n9854_o;
  wire n9855_o;
  wire n9856_o;
  wire n9857_o;
  wire n9858_o;
  wire n9859_o;
  wire n9860_o;
  wire n9861_o;
  wire n9862_o;
  wire n9863_o;
  wire n9864_o;
  wire n9865_o;
  wire n9866_o;
  wire n9867_o;
  wire n9868_o;
  wire n9869_o;
  wire n9870_o;
  wire n9871_o;
  wire n9872_o;
  wire n9873_o;
  wire n9874_o;
  wire n9875_o;
  wire n9876_o;
  wire n9877_o;
  wire n9878_o;
  wire n9879_o;
  wire n9880_o;
  wire n9881_o;
  wire n9882_o;
  wire n9883_o;
  wire n9884_o;
  wire n9885_o;
  wire n9886_o;
  wire [7:0] n9887_o;
  wire n9888_o;
  wire n9889_o;
  wire n9890_o;
  wire n9891_o;
  wire n9892_o;
  wire n9893_o;
  wire n9894_o;
  wire n9895_o;
  wire n9896_o;
  wire n9897_o;
  wire n9898_o;
  wire n9899_o;
  wire n9900_o;
  wire n9901_o;
  wire n9902_o;
  wire n9903_o;
  wire n9904_o;
  wire n9905_o;
  wire n9906_o;
  wire n9907_o;
  wire n9908_o;
  wire n9909_o;
  wire n9910_o;
  wire n9911_o;
  wire n9912_o;
  wire n9913_o;
  wire n9914_o;
  wire n9915_o;
  wire n9916_o;
  wire n9917_o;
  wire n9918_o;
  wire n9919_o;
  wire n9920_o;
  wire n9921_o;
  wire [7:0] n9922_o;
  wire n9923_o;
  wire n9924_o;
  wire n9925_o;
  wire n9926_o;
  wire n9927_o;
  wire n9928_o;
  wire n9929_o;
  wire n9930_o;
  wire n9931_o;
  wire n9932_o;
  wire n9933_o;
  wire n9934_o;
  wire n9935_o;
  wire n9936_o;
  wire n9937_o;
  wire n9938_o;
  wire n9939_o;
  wire n9940_o;
  wire n9941_o;
  wire n9942_o;
  wire n9943_o;
  wire n9944_o;
  wire n9945_o;
  wire n9946_o;
  wire n9947_o;
  wire n9948_o;
  wire n9949_o;
  wire n9950_o;
  wire n9951_o;
  wire n9952_o;
  wire n9953_o;
  wire n9954_o;
  wire n9955_o;
  wire n9956_o;
  wire [7:0] n9957_o;
  wire [6:0] n9958_o;
  wire n9959_o;
  wire n9960_o;
  wire n9961_o;
  wire n9962_o;
  wire n9963_o;
  wire n9964_o;
  wire n9965_o;
  wire n9966_o;
  wire n9967_o;
  wire n9968_o;
  wire n9969_o;
  wire n9970_o;
  wire n9971_o;
  wire n9972_o;
  wire n9973_o;
  wire n9974_o;
  wire n9975_o;
  wire n9976_o;
  wire n9977_o;
  wire n9978_o;
  wire n9979_o;
  wire n9980_o;
  wire n9981_o;
  wire n9982_o;
  wire n9983_o;
  wire n9984_o;
  wire n9985_o;
  wire n9986_o;
  wire n9987_o;
  wire n9988_o;
  wire n9989_o;
  wire n9990_o;
  wire n9991_o;
  wire n9992_o;
  wire n9993_o;
  wire n9994_o;
  wire n9995_o;
  wire n9996_o;
  wire n9997_o;
  wire n9998_o;
  wire n9999_o;
  wire n10000_o;
  wire n10001_o;
  wire n10002_o;
  wire n10003_o;
  wire n10004_o;
  wire n10005_o;
  wire n10006_o;
  wire n10007_o;
  wire n10008_o;
  wire n10009_o;
  wire n10010_o;
  wire n10011_o;
  wire n10012_o;
  wire n10013_o;
  wire n10014_o;
  wire n10015_o;
  wire n10016_o;
  wire n10017_o;
  wire n10018_o;
  wire n10019_o;
  wire n10020_o;
  wire n10021_o;
  wire n10022_o;
  wire n10023_o;
  wire n10024_o;
  wire n10025_o;
  wire n10026_o;
  wire n10027_o;
  wire n10028_o;
  wire n10029_o;
  wire n10030_o;
  wire n10031_o;
  wire n10032_o;
  wire n10033_o;
  wire n10034_o;
  wire n10035_o;
  wire n10036_o;
  wire n10037_o;
  wire n10038_o;
  wire n10039_o;
  wire n10040_o;
  wire n10041_o;
  wire n10042_o;
  wire n10043_o;
  wire n10044_o;
  wire n10045_o;
  wire n10046_o;
  wire n10047_o;
  wire n10048_o;
  wire n10049_o;
  wire n10050_o;
  wire n10051_o;
  wire n10052_o;
  wire n10053_o;
  wire n10054_o;
  wire n10055_o;
  wire n10056_o;
  wire n10057_o;
  wire n10058_o;
  wire n10059_o;
  wire n10060_o;
  wire n10061_o;
  wire n10062_o;
  wire n10063_o;
  wire n10064_o;
  wire n10065_o;
  wire n10066_o;
  wire n10067_o;
  wire n10068_o;
  wire n10069_o;
  wire n10070_o;
  wire n10071_o;
  wire n10072_o;
  wire n10073_o;
  wire n10074_o;
  wire n10075_o;
  wire n10076_o;
  wire n10077_o;
  wire n10078_o;
  wire n10079_o;
  wire n10080_o;
  wire n10081_o;
  wire n10082_o;
  wire n10083_o;
  wire n10084_o;
  wire n10085_o;
  wire n10086_o;
  wire n10087_o;
  wire n10088_o;
  wire n10089_o;
  wire n10090_o;
  wire n10091_o;
  wire n10092_o;
  wire n10093_o;
  wire n10094_o;
  wire n10095_o;
  wire n10096_o;
  wire n10097_o;
  wire n10098_o;
  wire n10099_o;
  wire n10100_o;
  wire n10101_o;
  wire n10102_o;
  wire n10103_o;
  wire n10104_o;
  wire n10105_o;
  wire n10106_o;
  wire n10107_o;
  wire n10108_o;
  wire n10109_o;
  wire n10110_o;
  wire n10111_o;
  wire n10112_o;
  wire n10113_o;
  wire n10114_o;
  wire n10115_o;
  wire n10116_o;
  wire n10117_o;
  wire n10118_o;
  wire n10119_o;
  wire n10120_o;
  wire n10121_o;
  wire n10122_o;
  wire n10123_o;
  wire n10124_o;
  wire n10125_o;
  wire n10126_o;
  wire n10127_o;
  wire n10128_o;
  wire n10129_o;
  wire n10130_o;
  wire n10131_o;
  wire n10132_o;
  wire n10133_o;
  wire n10134_o;
  wire n10135_o;
  wire n10136_o;
  wire n10137_o;
  wire n10138_o;
  wire n10139_o;
  wire n10140_o;
  wire n10141_o;
  wire n10142_o;
  wire n10143_o;
  wire n10144_o;
  wire n10145_o;
  wire n10146_o;
  wire n10147_o;
  wire n10148_o;
  wire n10149_o;
  wire n10150_o;
  wire n10151_o;
  wire n10152_o;
  wire n10153_o;
  wire n10154_o;
  wire n10155_o;
  wire n10156_o;
  wire n10157_o;
  wire n10158_o;
  wire n10159_o;
  wire n10160_o;
  wire n10161_o;
  wire n10162_o;
  wire n10163_o;
  wire n10164_o;
  wire n10165_o;
  wire n10166_o;
  wire n10167_o;
  wire n10168_o;
  wire n10169_o;
  wire n10170_o;
  wire n10171_o;
  wire n10172_o;
  wire n10173_o;
  wire n10174_o;
  wire n10175_o;
  wire n10176_o;
  wire n10177_o;
  wire n10178_o;
  wire n10179_o;
  wire n10180_o;
  wire n10181_o;
  wire n10182_o;
  wire n10183_o;
  wire n10184_o;
  wire n10185_o;
  wire n10186_o;
  wire n10187_o;
  wire n10188_o;
  wire n10189_o;
  wire n10190_o;
  wire n10191_o;
  wire n10192_o;
  wire n10193_o;
  wire n10194_o;
  wire n10195_o;
  wire n10196_o;
  wire n10197_o;
  wire n10198_o;
  wire n10199_o;
  wire n10200_o;
  wire n10201_o;
  wire n10202_o;
  wire n10203_o;
  wire n10204_o;
  wire n10205_o;
  wire n10206_o;
  wire n10207_o;
  wire n10208_o;
  wire n10209_o;
  wire n10210_o;
  wire n10211_o;
  wire n10212_o;
  wire n10213_o;
  wire n10214_o;
  wire n10215_o;
  wire n10216_o;
  wire n10217_o;
  wire n10218_o;
  wire n10219_o;
  wire n10220_o;
  wire n10221_o;
  wire n10222_o;
  wire n10223_o;
  wire n10224_o;
  wire n10225_o;
  wire n10226_o;
  wire n10227_o;
  wire n10228_o;
  wire n10229_o;
  wire n10230_o;
  wire n10231_o;
  wire n10232_o;
  wire n10233_o;
  wire n10234_o;
  wire n10235_o;
  wire n10236_o;
  wire n10237_o;
  wire n10238_o;
  wire n10239_o;
  wire n10240_o;
  wire n10241_o;
  wire n10242_o;
  wire n10243_o;
  wire n10244_o;
  wire n10245_o;
  wire n10246_o;
  wire n10247_o;
  wire n10248_o;
  wire n10249_o;
  wire n10250_o;
  wire n10251_o;
  wire n10252_o;
  wire n10253_o;
  wire n10254_o;
  wire n10255_o;
  wire n10256_o;
  wire n10257_o;
  wire n10258_o;
  wire n10259_o;
  wire n10260_o;
  wire n10261_o;
  wire n10262_o;
  wire n10263_o;
  wire n10264_o;
  wire n10265_o;
  wire n10266_o;
  wire n10267_o;
  wire n10268_o;
  wire n10269_o;
  wire n10270_o;
  wire n10271_o;
  wire n10272_o;
  wire n10273_o;
  wire n10274_o;
  wire n10275_o;
  wire n10276_o;
  wire n10277_o;
  wire n10278_o;
  wire n10279_o;
  wire n10280_o;
  wire n10281_o;
  wire n10282_o;
  wire n10283_o;
  wire n10284_o;
  wire n10285_o;
  wire n10286_o;
  wire n10287_o;
  wire n10288_o;
  wire n10289_o;
  wire n10290_o;
  wire n10291_o;
  wire n10292_o;
  wire n10293_o;
  wire n10294_o;
  wire n10295_o;
  wire n10296_o;
  wire n10297_o;
  wire n10298_o;
  wire n10299_o;
  wire n10300_o;
  wire n10301_o;
  wire n10302_o;
  wire n10303_o;
  wire n10304_o;
  wire n10305_o;
  wire n10306_o;
  wire n10307_o;
  wire n10308_o;
  wire n10309_o;
  wire n10310_o;
  wire n10311_o;
  wire n10312_o;
  wire n10313_o;
  wire n10314_o;
  wire n10315_o;
  wire n10316_o;
  wire n10317_o;
  wire n10318_o;
  wire n10319_o;
  wire n10320_o;
  wire n10321_o;
  wire n10322_o;
  wire n10323_o;
  wire n10324_o;
  wire n10325_o;
  wire n10326_o;
  wire n10327_o;
  wire n10328_o;
  wire n10329_o;
  wire n10330_o;
  wire n10331_o;
  wire n10332_o;
  wire n10333_o;
  wire n10334_o;
  wire n10335_o;
  wire n10336_o;
  wire n10337_o;
  wire n10338_o;
  wire n10339_o;
  wire n10340_o;
  wire n10341_o;
  wire n10342_o;
  wire n10343_o;
  wire n10344_o;
  wire n10345_o;
  wire n10346_o;
  wire n10347_o;
  wire n10348_o;
  wire n10349_o;
  wire n10350_o;
  wire n10351_o;
  wire n10352_o;
  wire n10353_o;
  wire n10354_o;
  wire n10355_o;
  wire n10356_o;
  wire n10357_o;
  wire n10358_o;
  wire n10359_o;
  wire n10360_o;
  wire n10361_o;
  wire n10362_o;
  wire n10363_o;
  wire n10364_o;
  wire n10365_o;
  wire n10366_o;
  wire n10367_o;
  wire n10368_o;
  wire n10369_o;
  wire n10370_o;
  wire n10371_o;
  wire n10372_o;
  wire n10373_o;
  wire n10374_o;
  wire n10375_o;
  wire n10376_o;
  wire n10377_o;
  wire n10378_o;
  wire n10379_o;
  wire n10380_o;
  wire n10381_o;
  wire n10382_o;
  wire n10383_o;
  wire n10384_o;
  wire n10385_o;
  wire n10386_o;
  wire n10387_o;
  wire n10388_o;
  wire n10389_o;
  wire n10390_o;
  wire n10391_o;
  wire n10392_o;
  wire n10393_o;
  wire n10394_o;
  wire n10395_o;
  wire n10396_o;
  wire n10397_o;
  wire n10398_o;
  wire n10399_o;
  wire n10400_o;
  wire n10401_o;
  wire n10402_o;
  wire n10403_o;
  wire n10404_o;
  wire n10405_o;
  wire n10406_o;
  wire n10407_o;
  wire n10408_o;
  wire n10409_o;
  wire n10410_o;
  wire n10411_o;
  wire n10412_o;
  wire n10413_o;
  wire n10414_o;
  wire n10415_o;
  wire n10416_o;
  wire n10417_o;
  wire n10418_o;
  wire n10419_o;
  wire n10420_o;
  wire n10421_o;
  wire n10422_o;
  wire n10423_o;
  wire n10424_o;
  wire n10425_o;
  wire n10426_o;
  wire n10427_o;
  wire n10428_o;
  wire n10429_o;
  wire n10430_o;
  wire n10431_o;
  wire n10432_o;
  wire n10433_o;
  wire n10434_o;
  wire n10435_o;
  wire n10436_o;
  wire n10437_o;
  wire n10438_o;
  wire n10439_o;
  wire n10440_o;
  wire n10441_o;
  wire n10442_o;
  wire n10443_o;
  wire n10444_o;
  wire n10445_o;
  wire n10446_o;
  wire n10447_o;
  wire n10448_o;
  wire n10449_o;
  wire n10450_o;
  wire n10451_o;
  wire n10452_o;
  wire n10453_o;
  wire n10454_o;
  wire n10455_o;
  wire n10456_o;
  wire n10457_o;
  wire n10458_o;
  wire n10459_o;
  wire n10460_o;
  wire n10461_o;
  wire n10462_o;
  wire n10463_o;
  wire n10464_o;
  wire n10465_o;
  wire n10466_o;
  wire n10467_o;
  wire n10468_o;
  wire n10469_o;
  wire n10470_o;
  wire n10471_o;
  wire n10472_o;
  wire n10473_o;
  wire n10474_o;
  wire n10475_o;
  wire n10476_o;
  wire n10477_o;
  wire n10478_o;
  wire n10479_o;
  wire n10480_o;
  wire [127:0] n10481_o;
  assign pc_o = pc_comb;
  assign ram_data_o = s_data;
  assign ram_adr_o = n7284_o;
  assign reg_data_o = s_reg_data;
  assign ram_wr_o = n8093_o;
  assign cy_o = n9136_o;
  assign ov_o = n7286_o;
  assign ram_en_o = n8928_o;
  assign acc_o = acc;
  assign p0_o = p0;
  assign p1_o = p1;
  assign p2_o = p2;
  assign p3_o = p3;
  assign all_trans_o = n9138_q;
  assign all_scon_o = n9139_o;
  assign all_sbuf_o = sbuf;
  assign all_smod_o = s_smodreg;
  assign all_tcon_tr0_o = n7302_o;
  assign all_tcon_tr1_o = n7303_o;
  assign all_tmod_o = tmod;
  assign all_reload_o = s_reload;
  assign all_wt_o = s_wt;
  assign all_wt_en_o = n9141_q;
  assign state_o = state;
  assign help_o = s_help;
  assign bit_data_o = s_bit_data;
  assign command_o = s_command;
  assign inthigh_o = s_inthigh;
  assign intlow_o = s_intlow;
  assign intpre_o = s_intpre;
  assign intpre2_o = s_intpre2;
  assign intblock_o = s_intblock_o;
  assign ti_o = s_ti;
  assign ri_o = s_ri;
  assign ie0_o = s_ie0;
  assign ie1_o = s_ie1;
  assign tf0_o = s_tf0;
  assign tf1_o = s_tf1;
  assign psw_o = psw;
  assign ie_o = ie;
  assign ip_o = ip;
  assign adrx_o = n9142_o;
  assign datax_o = acc;
  assign wrx_o = wrx_mux_i;
  assign memx_o = n8054_o;
  /* control_mem_rtl.vhd:74:11  */
  assign s_help = n8997_q; // (signal)
  /* control_mem_rtl.vhd:75:11  */
  assign s_help16 = n8999_q; // (signal)
  /* control_mem_rtl.vhd:76:11  */
  assign s_helpb = n9001_q; // (signal)
  /* control_mem_rtl.vhd:77:11  */
  assign s_ir = n9004_q; // (signal)
  /* control_mem_rtl.vhd:78:11  */
  assign gprbit = n9006_q; // (signal)
  /* control_mem_rtl.vhd:79:11  */
  assign s_r0_b0 = n9008_q; // (signal)
  /* control_mem_rtl.vhd:80:11  */
  assign s_r1_b0 = n9010_q; // (signal)
  /* control_mem_rtl.vhd:81:11  */
  assign s_r0_b1 = n9012_q; // (signal)
  /* control_mem_rtl.vhd:82:11  */
  assign s_r1_b1 = n9014_q; // (signal)
  /* control_mem_rtl.vhd:83:11  */
  assign s_r0_b2 = n9016_q; // (signal)
  /* control_mem_rtl.vhd:84:11  */
  assign s_r1_b2 = n9018_q; // (signal)
  /* control_mem_rtl.vhd:85:11  */
  assign s_r0_b3 = n9020_q; // (signal)
  /* control_mem_rtl.vhd:86:11  */
  assign s_r1_b3 = n9022_q; // (signal)
  /* control_mem_rtl.vhd:87:11  */
  assign s_reg_data = n7665_o; // (signal)
  /* control_mem_rtl.vhd:88:11  */
  assign state = n9024_q; // (signal)
  /* control_mem_rtl.vhd:340:50  */
  assign s_command = n7339_o; // (signal)
  /* control_mem_rtl.vhd:91:11  */
  assign s_pc_inc_en = pc_inc_en_i; // (signal)
  /* control_mem_rtl.vhd:92:11  */
  assign s_regs_wr_en = regs_wr_en_i; // (signal)
  /* control_mem_rtl.vhd:93:11  */
  assign s_data_mux = data_mux_i; // (signal)
  /* control_mem_rtl.vhd:94:11  */
  assign s_bdata_mux = bdata_mux_i; // (signal)
  /* control_mem_rtl.vhd:95:11  */
  assign s_adr_mux = adr_mux_i; // (signal)
  /* control_mem_rtl.vhd:96:11  */
  assign s_adrx_mux = adrx_mux_i; // (signal)
  /* control_mem_rtl.vhd:97:11  */
  assign s_help_en = help_en_i; // (signal)
  /* control_mem_rtl.vhd:98:11  */
  assign s_help16_en = help16_en_i; // (signal)
  /* control_mem_rtl.vhd:99:11  */
  assign s_helpb_en = helpb_en_i; // (signal)
  /* control_mem_rtl.vhd:100:11  */
  assign s_intpre2_d = intpre2_d_i; // (signal)
  /* control_mem_rtl.vhd:101:11  */
  assign s_intpre2_en = intpre2_en_i; // (signal)
  /* control_mem_rtl.vhd:102:11  */
  assign s_intlow_d = intlow_d_i; // (signal)
  /* control_mem_rtl.vhd:103:11  */
  assign s_intlow_en = intlow_en_i; // (signal)
  /* control_mem_rtl.vhd:104:11  */
  assign s_inthigh_d = inthigh_d_i; // (signal)
  /* control_mem_rtl.vhd:105:11  */
  assign s_inthigh_en = inthigh_en_i; // (signal)
  /* control_mem_rtl.vhd:106:11  */
  assign s_ext0isr_d = n9027_q; // (signal)
  /* control_mem_rtl.vhd:107:11  */
  assign s_ext0isrh_d = n9030_q; // (signal)
  /* control_mem_rtl.vhd:108:11  */
  assign s_ext1isr_d = n9033_q; // (signal)
  /* control_mem_rtl.vhd:109:11  */
  assign s_ext1isrh_d = n9036_q; // (signal)
  /* control_mem_rtl.vhd:111:11  */
  assign s_nextstate = nextstate_i; // (signal)
  /* control_mem_rtl.vhd:113:11  */
  assign s_bit_data = n7750_o; // (signal)
  /* control_mem_rtl.vhd:114:11  */
  assign s_intpre = n7877_o; // (signal)
  /* control_mem_rtl.vhd:115:11  */
  assign s_intpre2 = n9039_q; // (signal)
  /* control_mem_rtl.vhd:116:11  */
  assign s_inthigh = n9042_q; // (signal)
  /* control_mem_rtl.vhd:117:11  */
  assign s_intlow = n9045_q; // (signal)
  /* control_mem_rtl.vhd:118:11  */
  assign s_intblock = n7388_o; // (signal)
  /* control_mem_rtl.vhd:119:11  */
  assign s_intblock_o = n9047_q; // (signal)
  /* control_mem_rtl.vhd:959:67  */
  assign s_int0_edge = n7753_o; // (signal)
  /* control_mem_rtl.vhd:956:67  */
  assign s_int1_edge = n7755_o; // (signal)
  /* control_mem_rtl.vhd:962:49  */
  assign s_tf0_edge = n7757_o; // (signal)
  /* control_mem_rtl.vhd:963:49  */
  assign s_tf1_edge = n7759_o; // (signal)
  /* control_mem_rtl.vhd:967:48  */
  assign s_ri_edge = n7761_o; // (signal)
  /* control_mem_rtl.vhd:968:48  */
  assign s_ti_edge = n7763_o; // (signal)
  /* control_mem_rtl.vhd:322:21  */
  assign s_smodreg = n9049_q; // (signal)
  /* control_mem_rtl.vhd:415:47  */
  assign s_tl0 = all_tl0_i; // (signal)
  /* control_mem_rtl.vhd:416:47  */
  assign s_tl1 = all_tl1_i; // (signal)
  /* control_mem_rtl.vhd:417:47  */
  assign s_th0 = all_th0_i; // (signal)
  /* control_mem_rtl.vhd:418:47  */
  assign s_th1 = all_th1_i; // (signal)
  /* control_mem_rtl.vhd:430:49  */
  assign s_sbufi = all_sbuf_i; // (signal)
  /* control_mem_rtl.vhd:292:66  */
  assign s_reload = n9051_q; // (signal)
  /* control_mem_rtl.vhd:293:58  */
  assign s_wt = n9053_q; // (signal)
  /* control_mem_rtl.vhd:137:11  */
  assign s_tf1 = n7304_o; // (signal)
  /* control_mem_rtl.vhd:138:11  */
  assign s_tf0 = n7305_o; // (signal)
  /* control_mem_rtl.vhd:139:11  */
  assign s_ie1 = n7306_o; // (signal)
  /* control_mem_rtl.vhd:140:11  */
  assign s_ie0 = n7307_o; // (signal)
  /* control_mem_rtl.vhd:142:11  */
  assign s_ri = n7321_o; // (signal)
  /* control_mem_rtl.vhd:143:11  */
  assign s_ti = n7320_o; // (signal)
  /* control_mem_rtl.vhd:144:11  */
  assign s_rb8 = n7319_o; // (signal)
  /* control_mem_rtl.vhd:145:11  */
  assign s_tb8 = n7318_o; // (signal)
  /* control_mem_rtl.vhd:146:11  */
  assign s_ren = n7317_o; // (signal)
  /* control_mem_rtl.vhd:147:11  */
  assign s_sm2 = n7316_o; // (signal)
  /* control_mem_rtl.vhd:148:11  */
  assign s_sm1 = n7315_o; // (signal)
  /* control_mem_rtl.vhd:149:11  */
  assign s_sm0 = n7314_o; // (signal)
  /* control_mem_rtl.vhd:150:11  */
  assign s_smod = s_smodreg; // (signal)
  /* control_mem_rtl.vhd:558:34  */
  assign s_int0_h1 = n9055_q; // (signal)
  /* control_mem_rtl.vhd:960:59  */
  assign s_int0_h2 = n9057_q; // (signal)
  /* control_mem_rtl.vhd:500:53  */
  assign s_int0_h3 = n9059_q; // (signal)
  /* control_mem_rtl.vhd:561:34  */
  assign s_int1_h1 = n9061_q; // (signal)
  /* control_mem_rtl.vhd:957:59  */
  assign s_int1_h2 = n9063_q; // (signal)
  /* control_mem_rtl.vhd:502:53  */
  assign s_int1_h3 = n9065_q; // (signal)
  /* control_mem_rtl.vhd:566:32  */
  assign s_tf0_h1 = n9067_q; // (signal)
  /* control_mem_rtl.vhd:508:50  */
  assign s_tf0_h2 = n9069_q; // (signal)
  /* control_mem_rtl.vhd:568:32  */
  assign s_tf1_h1 = n9071_q; // (signal)
  /* control_mem_rtl.vhd:510:50  */
  assign s_tf1_h2 = n9073_q; // (signal)
  /* control_mem_rtl.vhd:573:30  */
  assign s_ri_h1 = n9075_q; // (signal)
  /* control_mem_rtl.vhd:516:47  */
  assign s_ri_h2 = n9077_q; // (signal)
  /* control_mem_rtl.vhd:575:30  */
  assign s_ti_h1 = n9079_q; // (signal)
  /* control_mem_rtl.vhd:518:47  */
  assign s_ti_h2 = n9081_q; // (signal)
  /* control_mem_rtl.vhd:167:11  */
  assign s_p = n7336_o; // (signal)
  /* control_mem_rtl.vhd:169:11  */
  assign s_p0 = n9085_q; // (signal)
  /* control_mem_rtl.vhd:170:11  */
  assign s_p1 = n9087_q; // (signal)
  /* control_mem_rtl.vhd:171:11  */
  assign s_p2 = n9089_q; // (signal)
  /* control_mem_rtl.vhd:172:11  */
  assign s_p3 = n9091_q; // (signal)
  /* control_mem_rtl.vhd:174:11  */
  assign pc = n9093_q; // (signal)
  /* control_mem_rtl.vhd:175:11  */
  assign pc_comb = n9094_o; // (signal)
  /* control_mem_rtl.vhd:176:11  */
  assign pc_plus1 = n7280_o; // (signal)
  /* control_mem_rtl.vhd:177:11  */
  assign pc_plus2 = n7283_o; // (signal)
  /* control_mem_rtl.vhd:179:11  */
  assign s_data = n9095_o; // (signal)
  /* control_mem_rtl.vhd:180:11  */
  assign s_adr = n8040_o; // (signal)
  /* control_mem_rtl.vhd:181:11  */
  assign s_preadr = n9097_q; // (signal)
  /* control_mem_rtl.vhd:182:11  */
  assign s_bdata = n7993_o; // (signal)
  /* control_mem_rtl.vhd:183:11  */
  assign s_rr_adr = n7344_o; // (signal)
  /* control_mem_rtl.vhd:184:11  */
  assign s_ri_adr = n7349_o; // (signal)
  /* control_mem_rtl.vhd:185:11  */
  assign s_ri_data = n8073_o; // (signal)
  /* control_mem_rtl.vhd:189:11  */
  assign p0 = n9099_q; // (signal)
  /* control_mem_rtl.vhd:190:11  */
  assign sp = n9101_q; // (signal)
  /* control_mem_rtl.vhd:191:11  */
  assign dpl = n9103_q; // (signal)
  /* control_mem_rtl.vhd:192:11  */
  assign dph = n9105_q; // (signal)
  /* control_mem_rtl.vhd:193:11  */
  assign pcon = n9107_q; // (signal)
  /* control_mem_rtl.vhd:413:55  */
  assign tcon = n9109_q; // (signal)
  /* control_mem_rtl.vhd:414:55  */
  assign tmod = n9111_q; // (signal)
  /* control_mem_rtl.vhd:196:11  */
  assign p1 = n9113_q; // (signal)
  /* control_mem_rtl.vhd:197:11  */
  assign scon = n9115_q; // (signal)
  /* control_mem_rtl.vhd:310:60  */
  assign sbuf = n9117_q; // (signal)
  /* control_mem_rtl.vhd:199:11  */
  assign p2 = n9119_q; // (signal)
  /* control_mem_rtl.vhd:200:11  */
  assign ie = n9121_q; // (signal)
  /* control_mem_rtl.vhd:201:11  */
  assign p3 = n9123_q; // (signal)
  /* control_mem_rtl.vhd:202:11  */
  assign ip = n9125_q; // (signal)
  /* control_mem_rtl.vhd:203:11  */
  assign psw = n9127_q; // (signal)
  /* control_mem_rtl.vhd:204:11  */
  assign acc = n9129_q; // (signal)
  /* control_mem_rtl.vhd:205:11  */
  assign b = n9131_q; // (signal)
  /* control_mem_rtl.vhd:209:11  */
  assign tsel = n9133_q; // (signal)
  /* control_mem_rtl.vhd:210:11  */
  assign ssel = n9135_q; // (signal)
  /* control_mem_rtl.vhd:232:18  */
  assign n7280_o = pc + 16'b0000000000000001;
  /* control_mem_rtl.vhd:233:18  */
  assign n7283_o = pc + 16'b0000000000000010;
  /* control_mem_rtl.vhd:234:38  */
  assign n7284_o = s_adr[6:0];
  assign n7285_o = psw[7];
  assign n7286_o = psw[2];
  assign n7287_o = psw[6];
  /* control_mem_rtl.vhd:285:33  */
  assign n7302_o = tcon[4];
  /* control_mem_rtl.vhd:286:33  */
  assign n7303_o = tcon[6];
  /* control_mem_rtl.vhd:296:24  */
  assign n7304_o = tcon[7];
  /* control_mem_rtl.vhd:297:24  */
  assign n7305_o = tcon[5];
  /* control_mem_rtl.vhd:298:24  */
  assign n7306_o = tcon[3];
  /* control_mem_rtl.vhd:299:24  */
  assign n7307_o = tcon[1];
  /* control_mem_rtl.vhd:303:35  */
  assign n7308_o = scon[0];
  /* control_mem_rtl.vhd:304:35  */
  assign n7309_o = scon[7];
  /* control_mem_rtl.vhd:305:35  */
  assign n7310_o = scon[6];
  /* control_mem_rtl.vhd:306:35  */
  assign n7311_o = scon[5];
  /* control_mem_rtl.vhd:307:35  */
  assign n7312_o = scon[4];
  /* control_mem_rtl.vhd:308:31  */
  assign n7313_o = scon[3];
  /* control_mem_rtl.vhd:314:24  */
  assign n7314_o = scon[7];
  /* control_mem_rtl.vhd:315:24  */
  assign n7315_o = scon[6];
  /* control_mem_rtl.vhd:316:24  */
  assign n7316_o = scon[5];
  /* control_mem_rtl.vhd:317:24  */
  assign n7317_o = scon[4];
  /* control_mem_rtl.vhd:318:24  */
  assign n7318_o = scon[3];
  /* control_mem_rtl.vhd:319:22  */
  assign n7319_o = all_scon_i[2];
  /* control_mem_rtl.vhd:320:24  */
  assign n7320_o = scon[1];
  /* control_mem_rtl.vhd:321:24  */
  assign n7321_o = scon[0];
  /* control_mem_rtl.vhd:329:13  */
  assign n7322_o = acc[7];
  /* control_mem_rtl.vhd:329:24  */
  assign n7323_o = acc[6];
  /* control_mem_rtl.vhd:329:17  */
  assign n7324_o = n7322_o ^ n7323_o;
  /* control_mem_rtl.vhd:329:35  */
  assign n7325_o = acc[5];
  /* control_mem_rtl.vhd:329:28  */
  assign n7326_o = n7324_o ^ n7325_o;
  /* control_mem_rtl.vhd:329:46  */
  assign n7327_o = acc[4];
  /* control_mem_rtl.vhd:329:39  */
  assign n7328_o = n7326_o ^ n7327_o;
  /* control_mem_rtl.vhd:330:13  */
  assign n7329_o = acc[3];
  /* control_mem_rtl.vhd:329:50  */
  assign n7330_o = n7328_o ^ n7329_o;
  /* control_mem_rtl.vhd:330:24  */
  assign n7331_o = acc[2];
  /* control_mem_rtl.vhd:330:17  */
  assign n7332_o = n7330_o ^ n7331_o;
  /* control_mem_rtl.vhd:330:35  */
  assign n7333_o = acc[1];
  /* control_mem_rtl.vhd:330:28  */
  assign n7334_o = n7332_o ^ n7333_o;
  /* control_mem_rtl.vhd:330:46  */
  assign n7335_o = acc[0];
  /* control_mem_rtl.vhd:330:39  */
  assign n7336_o = n7334_o ^ n7335_o;
  /* control_mem_rtl.vhd:334:37  */
  assign n7338_o = state == 3'b001;
  /* control_mem_rtl.vhd:334:27  */
  assign n7339_o = n7338_o ? rom_data_i : s_ir;
  /* control_mem_rtl.vhd:337:29  */
  assign n7341_o = psw & 8'b00011000;
  /* control_mem_rtl.vhd:338:15  */
  assign n7343_o = rom_data_i & 8'b00000111;
  /* control_mem_rtl.vhd:337:45  */
  assign n7344_o = n7341_o | n7343_o;
  /* control_mem_rtl.vhd:340:21  */
  assign n7346_o = psw & 8'b00011000;
  /* control_mem_rtl.vhd:340:63  */
  assign n7348_o = s_command & 8'b00000001;
  /* control_mem_rtl.vhd:340:37  */
  assign n7349_o = n7346_o | n7348_o;
  /* control_mem_rtl.vhd:368:41  */
  assign n7353_o = s_command == 8'b00110010;
  /* control_mem_rtl.vhd:370:27  */
  assign n7355_o = s_regs_wr_en == 3'b100;
  /* control_mem_rtl.vhd:371:14  */
  assign n7356_o = {24'b0, s_adr};  //  uext
  /* control_mem_rtl.vhd:371:34  */
  assign n7358_o = n7356_o == 32'b00000000000000000000000010111000;
  /* control_mem_rtl.vhd:371:46  */
  assign n7359_o = {24'b0, s_adr};  //  uext
  /* control_mem_rtl.vhd:371:66  */
  assign n7361_o = n7359_o == 32'b00000000000000000000000010101000;
  /* control_mem_rtl.vhd:371:43  */
  assign n7362_o = n7358_o | n7361_o;
  /* control_mem_rtl.vhd:370:35  */
  assign n7363_o = n7355_o & n7362_o;
  /* control_mem_rtl.vhd:372:24  */
  assign n7364_o = ~s_intpre2;
  /* control_mem_rtl.vhd:371:76  */
  assign n7365_o = n7363_o & n7364_o;
  /* control_mem_rtl.vhd:369:11  */
  assign n7366_o = n7353_o | n7365_o;
  /* control_mem_rtl.vhd:374:27  */
  assign n7368_o = s_regs_wr_en == 3'b110;
  /* control_mem_rtl.vhd:375:19  */
  assign n7369_o = s_adr[7:3];
  /* control_mem_rtl.vhd:375:32  */
  assign n7371_o = n7369_o == 5'b10101;
  /* control_mem_rtl.vhd:375:62  */
  assign n7372_o = s_adr[7:3];
  /* control_mem_rtl.vhd:375:75  */
  assign n7374_o = n7372_o == 5'b10111;
  /* control_mem_rtl.vhd:375:54  */
  assign n7375_o = n7371_o | n7374_o;
  /* control_mem_rtl.vhd:374:35  */
  assign n7376_o = n7368_o & n7375_o;
  /* control_mem_rtl.vhd:376:24  */
  assign n7377_o = ~s_intpre2;
  /* control_mem_rtl.vhd:375:98  */
  assign n7378_o = n7376_o & n7377_o;
  /* control_mem_rtl.vhd:373:11  */
  assign n7379_o = n7366_o | n7378_o;
  /* control_mem_rtl.vhd:379:28  */
  assign n7381_o = s_nextstate == 3'b001;
  /* control_mem_rtl.vhd:379:69  */
  assign n7383_o = s_command != 8'b00110010;
  /* control_mem_rtl.vhd:379:36  */
  assign n7384_o = n7381_o & n7383_o;
  /* control_mem_rtl.vhd:379:9  */
  assign n7386_o = n7384_o ? 1'b0 : s_intblock_o;
  /* control_mem_rtl.vhd:368:9  */
  assign n7388_o = n7379_o ? 1'b1 : n7386_o;
  /* control_mem_rtl.vhd:403:16  */
  assign n7391_o = s_preadr[7];
  /* control_mem_rtl.vhd:404:12  */
  assign n7392_o = {24'b0, s_preadr};  //  uext
  /* control_mem_rtl.vhd:405:13  */
  assign n7394_o = n7392_o == 32'b00000000000000000000000010000000;
  /* control_mem_rtl.vhd:406:13  */
  assign n7396_o = n7392_o == 32'b00000000000000000000000010000001;
  /* control_mem_rtl.vhd:407:13  */
  assign n7398_o = n7392_o == 32'b00000000000000000000000010000010;
  /* control_mem_rtl.vhd:408:13  */
  assign n7400_o = n7392_o == 32'b00000000000000000000000010000011;
  /* control_mem_rtl.vhd:409:13  */
  assign n7403_o = n7392_o == 32'b00000000000000000000000010000111;
  /* control_mem_rtl.vhd:413:13  */
  assign n7405_o = n7392_o == 32'b00000000000000000000000010001000;
  /* control_mem_rtl.vhd:414:13  */
  assign n7407_o = n7392_o == 32'b00000000000000000000000010001001;
  /* control_mem_rtl.vhd:415:13  */
  assign n7409_o = n7392_o == 32'b00000000000000000000000010001010;
  /* control_mem_rtl.vhd:416:13  */
  assign n7411_o = n7392_o == 32'b00000000000000000000000010001011;
  /* control_mem_rtl.vhd:417:13  */
  assign n7413_o = n7392_o == 32'b00000000000000000000000010001100;
  /* control_mem_rtl.vhd:418:13  */
  assign n7415_o = n7392_o == 32'b00000000000000000000000010001101;
  /* control_mem_rtl.vhd:419:13  */
  assign n7417_o = n7392_o == 32'b00000000000000000000000010001110;
  /* control_mem_rtl.vhd:420:13  */
  assign n7419_o = n7392_o == 32'b00000000000000000000000010010000;
  /* control_mem_rtl.vhd:421:13  */
  assign n7421_o = n7392_o == 32'b00000000000000000000000010011000;
  /* control_mem_rtl.vhd:430:13  */
  assign n7423_o = n7392_o == 32'b00000000000000000000000010011001;
  /* control_mem_rtl.vhd:431:13  */
  assign n7425_o = n7392_o == 32'b00000000000000000000000010011010;
  /* control_mem_rtl.vhd:432:13  */
  assign n7427_o = n7392_o == 32'b00000000000000000000000010100000;
  /* control_mem_rtl.vhd:433:13  */
  assign n7429_o = n7392_o == 32'b00000000000000000000000010101000;
  /* control_mem_rtl.vhd:434:13  */
  assign n7431_o = n7392_o == 32'b00000000000000000000000010110000;
  /* control_mem_rtl.vhd:435:13  */
  assign n7433_o = n7392_o == 32'b00000000000000000000000010111000;
  /* control_mem_rtl.vhd:436:13  */
  assign n7435_o = n7392_o == 32'b00000000000000000000000011010000;
  /* control_mem_rtl.vhd:437:13  */
  assign n7437_o = n7392_o == 32'b00000000000000000000000011100000;
  /* control_mem_rtl.vhd:438:13  */
  assign n7439_o = n7392_o == 32'b00000000000000000000000011110000;
  assign n7440_o = {n7439_o, n7437_o, n7435_o, n7433_o, n7431_o, n7429_o, n7427_o, n7425_o, n7423_o, n7421_o, n7419_o, n7417_o, n7415_o, n7413_o, n7411_o, n7409_o, n7407_o, n7405_o, n7403_o, n7400_o, n7398_o, n7396_o, n7394_o};
  assign n7441_o = s_p0[0];
  assign n7442_o = sp[0];
  assign n7443_o = dpl[0];
  assign n7444_o = dph[0];
  assign n7445_o = pcon[0];
  assign n7446_o = tcon[0];
  assign n7447_o = tmod[0];
  assign n7448_o = s_tl0[0];
  assign n7449_o = s_tl1[0];
  assign n7450_o = s_th0[0];
  assign n7451_o = s_th1[0];
  assign n7452_o = tsel[0];
  assign n7453_o = s_p1[0];
  assign n7454_o = s_sbufi[0];
  assign n7455_o = ssel[0];
  assign n7456_o = s_p2[0];
  assign n7457_o = ie[0];
  assign n7458_o = s_p3[0];
  assign n7459_o = ip[0];
  assign n7460_o = psw[0];
  assign n7461_o = acc[0];
  assign n7462_o = b[0];
  /* control_mem_rtl.vhd:404:7  */
  always @*
    case (n7440_o)
      23'b10000000000000000000000: n7464_o = n7462_o;
      23'b01000000000000000000000: n7464_o = n7461_o;
      23'b00100000000000000000000: n7464_o = n7460_o;
      23'b00010000000000000000000: n7464_o = n7459_o;
      23'b00001000000000000000000: n7464_o = n7458_o;
      23'b00000100000000000000000: n7464_o = n7457_o;
      23'b00000010000000000000000: n7464_o = n7456_o;
      23'b00000001000000000000000: n7464_o = n7455_o;
      23'b00000000100000000000000: n7464_o = n7454_o;
      23'b00000000010000000000000: n7464_o = s_ri;
      23'b00000000001000000000000: n7464_o = n7453_o;
      23'b00000000000100000000000: n7464_o = n7452_o;
      23'b00000000000010000000000: n7464_o = n7451_o;
      23'b00000000000001000000000: n7464_o = n7450_o;
      23'b00000000000000100000000: n7464_o = n7449_o;
      23'b00000000000000010000000: n7464_o = n7448_o;
      23'b00000000000000001000000: n7464_o = n7447_o;
      23'b00000000000000000100000: n7464_o = n7446_o;
      23'b00000000000000000010000: n7464_o = n7445_o;
      23'b00000000000000000001000: n7464_o = n7444_o;
      23'b00000000000000000000100: n7464_o = n7443_o;
      23'b00000000000000000000010: n7464_o = n7442_o;
      23'b00000000000000000000001: n7464_o = n7441_o;
      default: n7464_o = 1'b0;
    endcase
  assign n7465_o = s_p0[1];
  assign n7466_o = sp[1];
  assign n7467_o = dpl[1];
  assign n7468_o = dph[1];
  assign n7469_o = pcon[1];
  assign n7470_o = tcon[1];
  assign n7471_o = tmod[1];
  assign n7472_o = s_tl0[1];
  assign n7473_o = s_tl1[1];
  assign n7474_o = s_th0[1];
  assign n7475_o = s_th1[1];
  assign n7476_o = tsel[1];
  assign n7477_o = s_p1[1];
  assign n7478_o = s_sbufi[1];
  assign n7479_o = ssel[1];
  assign n7480_o = s_p2[1];
  assign n7481_o = ie[1];
  assign n7482_o = s_p3[1];
  assign n7483_o = ip[1];
  assign n7484_o = psw[1];
  assign n7485_o = acc[1];
  assign n7486_o = b[1];
  /* control_mem_rtl.vhd:404:7  */
  always @*
    case (n7440_o)
      23'b10000000000000000000000: n7488_o = n7486_o;
      23'b01000000000000000000000: n7488_o = n7485_o;
      23'b00100000000000000000000: n7488_o = n7484_o;
      23'b00010000000000000000000: n7488_o = n7483_o;
      23'b00001000000000000000000: n7488_o = n7482_o;
      23'b00000100000000000000000: n7488_o = n7481_o;
      23'b00000010000000000000000: n7488_o = n7480_o;
      23'b00000001000000000000000: n7488_o = n7479_o;
      23'b00000000100000000000000: n7488_o = n7478_o;
      23'b00000000010000000000000: n7488_o = s_ti;
      23'b00000000001000000000000: n7488_o = n7477_o;
      23'b00000000000100000000000: n7488_o = n7476_o;
      23'b00000000000010000000000: n7488_o = n7475_o;
      23'b00000000000001000000000: n7488_o = n7474_o;
      23'b00000000000000100000000: n7488_o = n7473_o;
      23'b00000000000000010000000: n7488_o = n7472_o;
      23'b00000000000000001000000: n7488_o = n7471_o;
      23'b00000000000000000100000: n7488_o = n7470_o;
      23'b00000000000000000010000: n7488_o = n7469_o;
      23'b00000000000000000001000: n7488_o = n7468_o;
      23'b00000000000000000000100: n7488_o = n7467_o;
      23'b00000000000000000000010: n7488_o = n7466_o;
      23'b00000000000000000000001: n7488_o = n7465_o;
      default: n7488_o = 1'b0;
    endcase
  assign n7489_o = s_p0[2];
  assign n7490_o = sp[2];
  assign n7491_o = dpl[2];
  assign n7492_o = dph[2];
  assign n7493_o = pcon[2];
  assign n7494_o = tcon[2];
  assign n7495_o = tmod[2];
  assign n7496_o = s_tl0[2];
  assign n7497_o = s_tl1[2];
  assign n7498_o = s_th0[2];
  assign n7499_o = s_th1[2];
  assign n7500_o = tsel[2];
  assign n7501_o = s_p1[2];
  assign n7502_o = s_sbufi[2];
  assign n7503_o = ssel[2];
  assign n7504_o = s_p2[2];
  assign n7505_o = ie[2];
  assign n7506_o = s_p3[2];
  assign n7507_o = ip[2];
  assign n7508_o = psw[2];
  assign n7509_o = acc[2];
  assign n7510_o = b[2];
  /* control_mem_rtl.vhd:404:7  */
  always @*
    case (n7440_o)
      23'b10000000000000000000000: n7512_o = n7510_o;
      23'b01000000000000000000000: n7512_o = n7509_o;
      23'b00100000000000000000000: n7512_o = n7508_o;
      23'b00010000000000000000000: n7512_o = n7507_o;
      23'b00001000000000000000000: n7512_o = n7506_o;
      23'b00000100000000000000000: n7512_o = n7505_o;
      23'b00000010000000000000000: n7512_o = n7504_o;
      23'b00000001000000000000000: n7512_o = n7503_o;
      23'b00000000100000000000000: n7512_o = n7502_o;
      23'b00000000010000000000000: n7512_o = s_rb8;
      23'b00000000001000000000000: n7512_o = n7501_o;
      23'b00000000000100000000000: n7512_o = n7500_o;
      23'b00000000000010000000000: n7512_o = n7499_o;
      23'b00000000000001000000000: n7512_o = n7498_o;
      23'b00000000000000100000000: n7512_o = n7497_o;
      23'b00000000000000010000000: n7512_o = n7496_o;
      23'b00000000000000001000000: n7512_o = n7495_o;
      23'b00000000000000000100000: n7512_o = n7494_o;
      23'b00000000000000000010000: n7512_o = n7493_o;
      23'b00000000000000000001000: n7512_o = n7492_o;
      23'b00000000000000000000100: n7512_o = n7491_o;
      23'b00000000000000000000010: n7512_o = n7490_o;
      23'b00000000000000000000001: n7512_o = n7489_o;
      default: n7512_o = 1'b0;
    endcase
  assign n7513_o = s_p0[3];
  assign n7514_o = sp[3];
  assign n7515_o = dpl[3];
  assign n7516_o = dph[3];
  assign n7517_o = pcon[3];
  assign n7518_o = tcon[3];
  assign n7519_o = tmod[3];
  assign n7520_o = s_tl0[3];
  assign n7521_o = s_tl1[3];
  assign n7522_o = s_th0[3];
  assign n7523_o = s_th1[3];
  assign n7524_o = tsel[3];
  assign n7525_o = s_p1[3];
  assign n7526_o = s_sbufi[3];
  assign n7527_o = ssel[3];
  assign n7528_o = s_p2[3];
  assign n7529_o = ie[3];
  assign n7530_o = s_p3[3];
  assign n7531_o = ip[3];
  assign n7532_o = psw[3];
  assign n7533_o = acc[3];
  assign n7534_o = b[3];
  /* control_mem_rtl.vhd:404:7  */
  always @*
    case (n7440_o)
      23'b10000000000000000000000: n7536_o = n7534_o;
      23'b01000000000000000000000: n7536_o = n7533_o;
      23'b00100000000000000000000: n7536_o = n7532_o;
      23'b00010000000000000000000: n7536_o = n7531_o;
      23'b00001000000000000000000: n7536_o = n7530_o;
      23'b00000100000000000000000: n7536_o = n7529_o;
      23'b00000010000000000000000: n7536_o = n7528_o;
      23'b00000001000000000000000: n7536_o = n7527_o;
      23'b00000000100000000000000: n7536_o = n7526_o;
      23'b00000000010000000000000: n7536_o = s_tb8;
      23'b00000000001000000000000: n7536_o = n7525_o;
      23'b00000000000100000000000: n7536_o = n7524_o;
      23'b00000000000010000000000: n7536_o = n7523_o;
      23'b00000000000001000000000: n7536_o = n7522_o;
      23'b00000000000000100000000: n7536_o = n7521_o;
      23'b00000000000000010000000: n7536_o = n7520_o;
      23'b00000000000000001000000: n7536_o = n7519_o;
      23'b00000000000000000100000: n7536_o = n7518_o;
      23'b00000000000000000010000: n7536_o = n7517_o;
      23'b00000000000000000001000: n7536_o = n7516_o;
      23'b00000000000000000000100: n7536_o = n7515_o;
      23'b00000000000000000000010: n7536_o = n7514_o;
      23'b00000000000000000000001: n7536_o = n7513_o;
      default: n7536_o = 1'b0;
    endcase
  assign n7537_o = s_p0[4];
  assign n7538_o = sp[4];
  assign n7539_o = dpl[4];
  assign n7540_o = dph[4];
  assign n7541_o = n7401_o[0];
  assign n7542_o = tcon[4];
  assign n7543_o = tmod[4];
  assign n7544_o = s_tl0[4];
  assign n7545_o = s_tl1[4];
  assign n7546_o = s_th0[4];
  assign n7547_o = s_th1[4];
  assign n7548_o = tsel[4];
  assign n7549_o = s_p1[4];
  assign n7550_o = s_sbufi[4];
  assign n7551_o = ssel[4];
  assign n7552_o = s_p2[4];
  assign n7553_o = ie[4];
  assign n7554_o = s_p3[4];
  assign n7555_o = ip[4];
  assign n7556_o = psw[4];
  assign n7557_o = acc[4];
  assign n7558_o = b[4];
  /* control_mem_rtl.vhd:404:7  */
  always @*
    case (n7440_o)
      23'b10000000000000000000000: n7560_o = n7558_o;
      23'b01000000000000000000000: n7560_o = n7557_o;
      23'b00100000000000000000000: n7560_o = n7556_o;
      23'b00010000000000000000000: n7560_o = n7555_o;
      23'b00001000000000000000000: n7560_o = n7554_o;
      23'b00000100000000000000000: n7560_o = n7553_o;
      23'b00000010000000000000000: n7560_o = n7552_o;
      23'b00000001000000000000000: n7560_o = n7551_o;
      23'b00000000100000000000000: n7560_o = n7550_o;
      23'b00000000010000000000000: n7560_o = s_ren;
      23'b00000000001000000000000: n7560_o = n7549_o;
      23'b00000000000100000000000: n7560_o = n7548_o;
      23'b00000000000010000000000: n7560_o = n7547_o;
      23'b00000000000001000000000: n7560_o = n7546_o;
      23'b00000000000000100000000: n7560_o = n7545_o;
      23'b00000000000000010000000: n7560_o = n7544_o;
      23'b00000000000000001000000: n7560_o = n7543_o;
      23'b00000000000000000100000: n7560_o = n7542_o;
      23'b00000000000000000010000: n7560_o = n7541_o;
      23'b00000000000000000001000: n7560_o = n7540_o;
      23'b00000000000000000000100: n7560_o = n7539_o;
      23'b00000000000000000000010: n7560_o = n7538_o;
      23'b00000000000000000000001: n7560_o = n7537_o;
      default: n7560_o = 1'b0;
    endcase
  assign n7561_o = s_p0[5];
  assign n7562_o = sp[5];
  assign n7563_o = dpl[5];
  assign n7564_o = dph[5];
  assign n7565_o = n7401_o[1];
  assign n7566_o = tcon[5];
  assign n7567_o = tmod[5];
  assign n7568_o = s_tl0[5];
  assign n7569_o = s_tl1[5];
  assign n7570_o = s_th0[5];
  assign n7571_o = s_th1[5];
  assign n7572_o = tsel[5];
  assign n7573_o = s_p1[5];
  assign n7574_o = s_sbufi[5];
  assign n7575_o = ssel[5];
  assign n7576_o = s_p2[5];
  assign n7577_o = ie[5];
  assign n7578_o = s_p3[5];
  assign n7579_o = ip[5];
  assign n7580_o = psw[5];
  assign n7581_o = acc[5];
  assign n7582_o = b[5];
  /* control_mem_rtl.vhd:404:7  */
  always @*
    case (n7440_o)
      23'b10000000000000000000000: n7584_o = n7582_o;
      23'b01000000000000000000000: n7584_o = n7581_o;
      23'b00100000000000000000000: n7584_o = n7580_o;
      23'b00010000000000000000000: n7584_o = n7579_o;
      23'b00001000000000000000000: n7584_o = n7578_o;
      23'b00000100000000000000000: n7584_o = n7577_o;
      23'b00000010000000000000000: n7584_o = n7576_o;
      23'b00000001000000000000000: n7584_o = n7575_o;
      23'b00000000100000000000000: n7584_o = n7574_o;
      23'b00000000010000000000000: n7584_o = s_sm2;
      23'b00000000001000000000000: n7584_o = n7573_o;
      23'b00000000000100000000000: n7584_o = n7572_o;
      23'b00000000000010000000000: n7584_o = n7571_o;
      23'b00000000000001000000000: n7584_o = n7570_o;
      23'b00000000000000100000000: n7584_o = n7569_o;
      23'b00000000000000010000000: n7584_o = n7568_o;
      23'b00000000000000001000000: n7584_o = n7567_o;
      23'b00000000000000000100000: n7584_o = n7566_o;
      23'b00000000000000000010000: n7584_o = n7565_o;
      23'b00000000000000000001000: n7584_o = n7564_o;
      23'b00000000000000000000100: n7584_o = n7563_o;
      23'b00000000000000000000010: n7584_o = n7562_o;
      23'b00000000000000000000001: n7584_o = n7561_o;
      default: n7584_o = 1'b0;
    endcase
  assign n7585_o = s_p0[6];
  assign n7586_o = sp[6];
  assign n7587_o = dpl[6];
  assign n7588_o = dph[6];
  assign n7589_o = n7401_o[2];
  assign n7590_o = tcon[6];
  assign n7591_o = tmod[6];
  assign n7592_o = s_tl0[6];
  assign n7593_o = s_tl1[6];
  assign n7594_o = s_th0[6];
  assign n7595_o = s_th1[6];
  assign n7596_o = tsel[6];
  assign n7597_o = s_p1[6];
  assign n7598_o = s_sbufi[6];
  assign n7599_o = ssel[6];
  assign n7600_o = s_p2[6];
  assign n7601_o = ie[6];
  assign n7602_o = s_p3[6];
  assign n7603_o = ip[6];
  assign n7604_o = psw[6];
  assign n7605_o = acc[6];
  assign n7606_o = b[6];
  /* control_mem_rtl.vhd:404:7  */
  always @*
    case (n7440_o)
      23'b10000000000000000000000: n7608_o = n7606_o;
      23'b01000000000000000000000: n7608_o = n7605_o;
      23'b00100000000000000000000: n7608_o = n7604_o;
      23'b00010000000000000000000: n7608_o = n7603_o;
      23'b00001000000000000000000: n7608_o = n7602_o;
      23'b00000100000000000000000: n7608_o = n7601_o;
      23'b00000010000000000000000: n7608_o = n7600_o;
      23'b00000001000000000000000: n7608_o = n7599_o;
      23'b00000000100000000000000: n7608_o = n7598_o;
      23'b00000000010000000000000: n7608_o = s_sm1;
      23'b00000000001000000000000: n7608_o = n7597_o;
      23'b00000000000100000000000: n7608_o = n7596_o;
      23'b00000000000010000000000: n7608_o = n7595_o;
      23'b00000000000001000000000: n7608_o = n7594_o;
      23'b00000000000000100000000: n7608_o = n7593_o;
      23'b00000000000000010000000: n7608_o = n7592_o;
      23'b00000000000000001000000: n7608_o = n7591_o;
      23'b00000000000000000100000: n7608_o = n7590_o;
      23'b00000000000000000010000: n7608_o = n7589_o;
      23'b00000000000000000001000: n7608_o = n7588_o;
      23'b00000000000000000000100: n7608_o = n7587_o;
      23'b00000000000000000000010: n7608_o = n7586_o;
      23'b00000000000000000000001: n7608_o = n7585_o;
      default: n7608_o = 1'b0;
    endcase
  assign n7609_o = s_p0[7];
  assign n7610_o = sp[7];
  assign n7611_o = dpl[7];
  assign n7612_o = dph[7];
  assign n7613_o = tcon[7];
  assign n7614_o = tmod[7];
  assign n7615_o = s_tl0[7];
  assign n7616_o = s_tl1[7];
  assign n7617_o = s_th0[7];
  assign n7618_o = s_th1[7];
  assign n7619_o = tsel[7];
  assign n7620_o = s_p1[7];
  assign n7621_o = s_sbufi[7];
  assign n7622_o = ssel[7];
  assign n7623_o = s_p2[7];
  assign n7624_o = ie[7];
  assign n7625_o = s_p3[7];
  assign n7626_o = ip[7];
  assign n7627_o = psw[7];
  assign n7628_o = acc[7];
  assign n7629_o = b[7];
  /* control_mem_rtl.vhd:404:7  */
  always @*
    case (n7440_o)
      23'b10000000000000000000000: n7631_o = n7629_o;
      23'b01000000000000000000000: n7631_o = n7628_o;
      23'b00100000000000000000000: n7631_o = n7627_o;
      23'b00010000000000000000000: n7631_o = n7626_o;
      23'b00001000000000000000000: n7631_o = n7625_o;
      23'b00000100000000000000000: n7631_o = n7624_o;
      23'b00000010000000000000000: n7631_o = n7623_o;
      23'b00000001000000000000000: n7631_o = n7622_o;
      23'b00000000100000000000000: n7631_o = n7621_o;
      23'b00000000010000000000000: n7631_o = s_sm0;
      23'b00000000001000000000000: n7631_o = n7620_o;
      23'b00000000000100000000000: n7631_o = n7619_o;
      23'b00000000000010000000000: n7631_o = n7618_o;
      23'b00000000000001000000000: n7631_o = n7617_o;
      23'b00000000000000100000000: n7631_o = n7616_o;
      23'b00000000000000010000000: n7631_o = n7615_o;
      23'b00000000000000001000000: n7631_o = n7614_o;
      23'b00000000000000000100000: n7631_o = n7613_o;
      23'b00000000000000000010000: n7631_o = s_smod;
      23'b00000000000000000001000: n7631_o = n7612_o;
      23'b00000000000000000000100: n7631_o = n7611_o;
      23'b00000000000000000000010: n7631_o = n7610_o;
      23'b00000000000000000000001: n7631_o = n7609_o;
      default: n7631_o = 1'b0;
    endcase
  /* control_mem_rtl.vhd:442:41  */
  assign n7632_o = s_preadr[7:4];
  /* control_mem_rtl.vhd:442:56  */
  assign n7634_o = n7632_o == 4'b0010;
  /* control_mem_rtl.vhd:443:55  */
  assign n7635_o = s_preadr[3:0];
  /* control_mem_rtl.vhd:445:44  */
  assign n7640_o = s_preadr == 8'b00000000;
  /* control_mem_rtl.vhd:447:44  */
  assign n7642_o = s_preadr == 8'b00000001;
  /* control_mem_rtl.vhd:449:44  */
  assign n7644_o = s_preadr == 8'b00001000;
  /* control_mem_rtl.vhd:451:44  */
  assign n7646_o = s_preadr == 8'b00001001;
  /* control_mem_rtl.vhd:453:44  */
  assign n7648_o = s_preadr == 8'b00010000;
  /* control_mem_rtl.vhd:455:44  */
  assign n7650_o = s_preadr == 8'b00010001;
  /* control_mem_rtl.vhd:457:44  */
  assign n7652_o = s_preadr == 8'b00011000;
  /* control_mem_rtl.vhd:459:44  */
  assign n7654_o = s_preadr == 8'b00011001;
  /* control_mem_rtl.vhd:459:5  */
  assign n7655_o = n7654_o ? s_r1_b3 : ram_data_i;
  /* control_mem_rtl.vhd:457:5  */
  assign n7656_o = n7652_o ? s_r0_b3 : n7655_o;
  /* control_mem_rtl.vhd:455:5  */
  assign n7657_o = n7650_o ? s_r1_b2 : n7656_o;
  /* control_mem_rtl.vhd:453:5  */
  assign n7658_o = n7648_o ? s_r0_b2 : n7657_o;
  /* control_mem_rtl.vhd:451:5  */
  assign n7659_o = n7646_o ? s_r1_b1 : n7658_o;
  /* control_mem_rtl.vhd:449:5  */
  assign n7660_o = n7644_o ? s_r0_b1 : n7659_o;
  /* control_mem_rtl.vhd:447:5  */
  assign n7661_o = n7642_o ? s_r1_b0 : n7660_o;
  /* control_mem_rtl.vhd:445:5  */
  assign n7662_o = n7640_o ? s_r0_b0 : n7661_o;
  /* control_mem_rtl.vhd:442:5  */
  assign n7663_o = n7634_o ? n9169_o : n7662_o;
  assign n7664_o = {n7631_o, n7608_o, n7584_o, n7560_o, n7536_o, n7512_o, n7488_o, n7464_o};
  /* control_mem_rtl.vhd:403:5  */
  assign n7665_o = n7391_o ? n7664_o : n7663_o;
  /* control_mem_rtl.vhd:466:16  */
  assign n7666_o = s_preadr[7];
  /* control_mem_rtl.vhd:467:20  */
  assign n7667_o = s_preadr[6:3];
  /* control_mem_rtl.vhd:468:64  */
  assign n7668_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:468:9  */
  assign n7673_o = n7667_o == 4'b0000;
  /* control_mem_rtl.vhd:470:59  */
  assign n7674_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:469:9  */
  assign n7679_o = n7667_o == 4'b0001;
  /* control_mem_rtl.vhd:471:64  */
  assign n7680_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:471:9  */
  assign n7685_o = n7667_o == 4'b0010;
  /* control_mem_rtl.vhd:473:35  */
  assign n7686_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:473:14  */
  assign n7687_o = {29'b0, n7686_o};  //  uext
  /* control_mem_rtl.vhd:473:48  */
  assign n7689_o = n7687_o == 32'b00000000000000000000000000000010;
  /* control_mem_rtl.vhd:476:61  */
  assign n7690_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:473:11  */
  assign n7694_o = n7689_o ? s_rb8 : n9225_o;
  /* control_mem_rtl.vhd:472:9  */
  assign n7696_o = n7667_o == 4'b0011;
  /* control_mem_rtl.vhd:478:64  */
  assign n7697_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:478:9  */
  assign n7702_o = n7667_o == 4'b0100;
  /* control_mem_rtl.vhd:479:62  */
  assign n7703_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:479:9  */
  assign n7708_o = n7667_o == 4'b0101;
  /* control_mem_rtl.vhd:480:64  */
  assign n7709_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:480:9  */
  assign n7714_o = n7667_o == 4'b0110;
  /* control_mem_rtl.vhd:481:62  */
  assign n7715_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:481:9  */
  assign n7720_o = n7667_o == 4'b0111;
  /* control_mem_rtl.vhd:482:63  */
  assign n7721_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:482:9  */
  assign n7726_o = n7667_o == 4'b1010;
  /* control_mem_rtl.vhd:483:63  */
  assign n7727_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:483:9  */
  assign n7732_o = n7667_o == 4'b1100;
  /* control_mem_rtl.vhd:484:61  */
  assign n7733_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:484:9  */
  assign n7738_o = n7667_o == 4'b1110;
  assign n7739_o = {n7738_o, n7732_o, n7726_o, n7720_o, n7714_o, n7708_o, n7702_o, n7696_o, n7685_o, n7679_o, n7673_o};
  /* control_mem_rtl.vhd:467:7  */
  always @*
    case (n7739_o)
      11'b10000000000: n7741_o = n9323_o;
      11'b01000000000: n7741_o = n9309_o;
      11'b00100000000: n7741_o = n9295_o;
      11'b00010000000: n7741_o = n9281_o;
      11'b00001000000: n7741_o = n9267_o;
      11'b00000100000: n7741_o = n9253_o;
      11'b00000010000: n7741_o = n9239_o;
      11'b00000001000: n7741_o = n7694_o;
      11'b00000000100: n7741_o = n9211_o;
      11'b00000000010: n7741_o = n9197_o;
      11'b00000000001: n7741_o = n9183_o;
      default: n7741_o = 1'b0;
    endcase
  /* control_mem_rtl.vhd:488:55  */
  assign n7742_o = s_preadr[6:3];
  /* control_mem_rtl.vhd:489:49  */
  assign n7745_o = s_preadr[2:0];
  /* control_mem_rtl.vhd:466:5  */
  assign n7750_o = n7666_o ? n7741_o : n9538_o;
  /* control_mem_rtl.vhd:500:23  */
  assign n7752_o = ~s_int0_h2;
  /* control_mem_rtl.vhd:500:40  */
  assign n7753_o = n7752_o & s_int0_h3;
  /* control_mem_rtl.vhd:502:23  */
  assign n7754_o = ~s_int1_h2;
  /* control_mem_rtl.vhd:502:40  */
  assign n7755_o = n7754_o & s_int1_h3;
  /* control_mem_rtl.vhd:508:38  */
  assign n7756_o = ~s_tf0_h2;
  /* control_mem_rtl.vhd:508:34  */
  assign n7757_o = s_tf0_h1 & n7756_o;
  /* control_mem_rtl.vhd:510:38  */
  assign n7758_o = ~s_tf1_h2;
  /* control_mem_rtl.vhd:510:34  */
  assign n7759_o = s_tf1_h1 & n7758_o;
  /* control_mem_rtl.vhd:516:36  */
  assign n7760_o = ~s_ri_h2;
  /* control_mem_rtl.vhd:516:32  */
  assign n7761_o = s_ri_h1 & n7760_o;
  /* control_mem_rtl.vhd:518:36  */
  assign n7762_o = ~s_ti_h2;
  /* control_mem_rtl.vhd:518:32  */
  assign n7763_o = s_ti_h1 & n7762_o;
  /* control_mem_rtl.vhd:572:33  */
  assign n7767_o = all_scon_i[0];
  /* control_mem_rtl.vhd:574:33  */
  assign n7768_o = all_scon_i[1];
  assign n7816_o = ie[7];
  assign n7817_o = ie[0];
  assign n7818_o = ie[1];
  /* control_mem_rtl.vhd:591:29  */
  assign n7819_o = n7817_o | n7818_o;
  assign n7820_o = ie[2];
  /* control_mem_rtl.vhd:591:40  */
  assign n7821_o = n7819_o | n7820_o;
  assign n7822_o = ie[3];
  /* control_mem_rtl.vhd:591:51  */
  assign n7823_o = n7821_o | n7822_o;
  assign n7824_o = ie[4];
  /* control_mem_rtl.vhd:591:62  */
  assign n7825_o = n7823_o | n7824_o;
  /* control_mem_rtl.vhd:591:16  */
  assign n7826_o = n7816_o & n7825_o;
  assign n7827_o = ie[0];
  assign n7828_o = ip[0];
  /* control_mem_rtl.vhd:595:18  */
  assign n7829_o = n7828_o & n7827_o;
  /* control_mem_rtl.vhd:595:26  */
  assign n7830_o = n7829_o & s_ie0;
  assign n7831_o = ie[1];
  assign n7832_o = ip[1];
  /* control_mem_rtl.vhd:596:18  */
  assign n7833_o = n7832_o & n7831_o;
  /* control_mem_rtl.vhd:596:26  */
  assign n7834_o = n7833_o & s_tf0;
  /* control_mem_rtl.vhd:595:37  */
  assign n7835_o = n7830_o | n7834_o;
  assign n7836_o = ie[2];
  assign n7837_o = ip[2];
  /* control_mem_rtl.vhd:597:18  */
  assign n7838_o = n7837_o & n7836_o;
  /* control_mem_rtl.vhd:597:26  */
  assign n7839_o = n7838_o & s_ie1;
  /* control_mem_rtl.vhd:596:37  */
  assign n7840_o = n7835_o | n7839_o;
  assign n7841_o = ie[3];
  assign n7842_o = ip[3];
  /* control_mem_rtl.vhd:598:18  */
  assign n7843_o = n7842_o & n7841_o;
  /* control_mem_rtl.vhd:598:26  */
  assign n7844_o = n7843_o & s_tf1;
  /* control_mem_rtl.vhd:597:37  */
  assign n7845_o = n7840_o | n7844_o;
  assign n7846_o = ie[4];
  assign n7847_o = ip[4];
  /* control_mem_rtl.vhd:599:18  */
  assign n7848_o = n7847_o & n7846_o;
  /* control_mem_rtl.vhd:599:35  */
  assign n7849_o = s_ri | s_ti;
  /* control_mem_rtl.vhd:599:25  */
  assign n7850_o = n7848_o & n7849_o;
  /* control_mem_rtl.vhd:598:37  */
  assign n7851_o = n7845_o | n7850_o;
  /* control_mem_rtl.vhd:595:9  */
  assign n7854_o = n7851_o ? 1'b1 : 1'b0;
  assign n7855_o = ie[0];
  /* control_mem_rtl.vhd:605:18  */
  assign n7856_o = n7855_o & s_ie0;
  assign n7857_o = ie[1];
  /* control_mem_rtl.vhd:606:18  */
  assign n7858_o = n7857_o & s_tf0;
  /* control_mem_rtl.vhd:605:29  */
  assign n7859_o = n7856_o | n7858_o;
  assign n7860_o = ie[2];
  /* control_mem_rtl.vhd:607:18  */
  assign n7861_o = n7860_o & s_ie1;
  /* control_mem_rtl.vhd:606:29  */
  assign n7862_o = n7859_o | n7861_o;
  assign n7863_o = ie[3];
  /* control_mem_rtl.vhd:608:18  */
  assign n7864_o = n7863_o & s_tf1;
  /* control_mem_rtl.vhd:607:29  */
  assign n7865_o = n7862_o | n7864_o;
  /* control_mem_rtl.vhd:609:27  */
  assign n7866_o = s_ri | s_ti;
  assign n7867_o = ie[4];
  /* control_mem_rtl.vhd:609:17  */
  assign n7868_o = n7867_o & n7866_o;
  /* control_mem_rtl.vhd:608:29  */
  assign n7869_o = n7865_o | n7868_o;
  /* control_mem_rtl.vhd:605:9  */
  assign n7872_o = n7869_o ? 1'b1 : 1'b0;
  /* control_mem_rtl.vhd:594:7  */
  assign n7873_o = s_intlow ? n7854_o : n7872_o;
  /* control_mem_rtl.vhd:592:7  */
  assign n7875_o = s_inthigh ? 1'b0 : n7873_o;
  /* control_mem_rtl.vhd:591:5  */
  assign n7877_o = n7826_o ? n7875_o : 1'b0;
  /* control_mem_rtl.vhd:638:7  */
  assign n7881_o = s_data_mux == 4'b0000;
  /* control_mem_rtl.vhd:639:34  */
  assign n7882_o = pc[7:0];
  /* control_mem_rtl.vhd:639:7  */
  assign n7884_o = s_data_mux == 4'b0001;
  /* control_mem_rtl.vhd:640:34  */
  assign n7885_o = pc[15:8];
  /* control_mem_rtl.vhd:640:7  */
  assign n7887_o = s_data_mux == 4'b0010;
  /* control_mem_rtl.vhd:641:7  */
  assign n7889_o = s_data_mux == 4'b0011;
  /* control_mem_rtl.vhd:642:7  */
  assign n7891_o = s_data_mux == 4'b0100;
  /* control_mem_rtl.vhd:643:7  */
  assign n7893_o = s_data_mux == 4'b0101;
  /* control_mem_rtl.vhd:644:7  */
  assign n7895_o = s_data_mux == 4'b0110;
  /* control_mem_rtl.vhd:646:34  */
  assign n7896_o = acc[3:0];
  /* control_mem_rtl.vhd:647:34  */
  assign n7897_o = acc[7:4];
  /* control_mem_rtl.vhd:645:7  */
  assign n7899_o = s_data_mux == 4'b0111;
  /* control_mem_rtl.vhd:648:7  */
  assign n7901_o = s_data_mux == 4'b1000;
  /* control_mem_rtl.vhd:650:41  */
  assign n7902_o = s_reg_data[7:4];
  /* control_mem_rtl.vhd:651:37  */
  assign n7903_o = s_help[3:0];
  /* control_mem_rtl.vhd:649:7  */
  assign n7905_o = s_data_mux == 4'b1001;
  /* control_mem_rtl.vhd:653:34  */
  assign n7906_o = acc[7:4];
  /* control_mem_rtl.vhd:654:41  */
  assign n7907_o = s_reg_data[3:0];
  /* control_mem_rtl.vhd:652:7  */
  assign n7909_o = s_data_mux == 4'b1010;
  /* control_mem_rtl.vhd:655:40  */
  assign n7910_o = s_help16[7:0];
  /* control_mem_rtl.vhd:655:7  */
  assign n7912_o = s_data_mux == 4'b1100;
  /* control_mem_rtl.vhd:656:40  */
  assign n7913_o = s_help16[15:8];
  /* control_mem_rtl.vhd:656:7  */
  assign n7915_o = s_data_mux == 4'b1101;
  /* control_mem_rtl.vhd:657:40  */
  assign n7916_o = pc_plus2[7:0];
  /* control_mem_rtl.vhd:657:7  */
  assign n7918_o = s_data_mux == 4'b1110;
  /* control_mem_rtl.vhd:658:7  */
  assign n7920_o = s_data_mux == 4'b1111;
  assign n7921_o = {n7920_o, n7918_o, n7915_o, n7912_o, n7909_o, n7905_o, n7901_o, n7899_o, n7895_o, n7893_o, n7891_o, n7889_o, n7887_o, n7884_o, n7881_o};
  assign n7923_o = n7882_o[3:0];
  assign n7924_o = n7885_o[3:0];
  assign n7925_o = aludata_i[3:0];
  assign n7926_o = s_reg_data[3:0];
  assign n7927_o = rom_data_i[3:0];
  assign n7928_o = acc[3:0];
  assign n7929_o = s_help[3:0];
  assign n7930_o = n7910_o[3:0];
  assign n7931_o = n7913_o[3:0];
  assign n7932_o = n7916_o[3:0];
  assign n7933_o = datax_i[3:0];
  /* control_mem_rtl.vhd:637:5  */
  always @*
    case (n7921_o)
      15'b100000000000000: n7935_o = n7933_o;
      15'b010000000000000: n7935_o = n7932_o;
      15'b001000000000000: n7935_o = n7931_o;
      15'b000100000000000: n7935_o = n7930_o;
      15'b000010000000000: n7935_o = n7907_o;
      15'b000001000000000: n7935_o = n7903_o;
      15'b000000100000000: n7935_o = n7929_o;
      15'b000000010000000: n7935_o = n7897_o;
      15'b000000001000000: n7935_o = n7928_o;
      15'b000000000100000: n7935_o = n7927_o;
      15'b000000000010000: n7935_o = n7926_o;
      15'b000000000001000: n7935_o = n7925_o;
      15'b000000000000100: n7935_o = n7924_o;
      15'b000000000000010: n7935_o = n7923_o;
      15'b000000000000001: n7935_o = 4'b0000;
      default: n7935_o = 4'b0000;
    endcase
  assign n7937_o = n7882_o[7:4];
  assign n7938_o = n7885_o[7:4];
  assign n7939_o = aludata_i[7:4];
  assign n7940_o = s_reg_data[7:4];
  assign n7941_o = rom_data_i[7:4];
  assign n7942_o = acc[7:4];
  assign n7943_o = s_help[7:4];
  assign n7944_o = n7910_o[7:4];
  assign n7945_o = n7913_o[7:4];
  assign n7946_o = n7916_o[7:4];
  assign n7947_o = datax_i[7:4];
  /* control_mem_rtl.vhd:637:5  */
  always @*
    case (n7921_o)
      15'b100000000000000: n7949_o = n7947_o;
      15'b010000000000000: n7949_o = n7946_o;
      15'b001000000000000: n7949_o = n7945_o;
      15'b000100000000000: n7949_o = n7944_o;
      15'b000010000000000: n7949_o = n7906_o;
      15'b000001000000000: n7949_o = n7902_o;
      15'b000000100000000: n7949_o = n7943_o;
      15'b000000010000000: n7949_o = n7896_o;
      15'b000000001000000: n7949_o = n7942_o;
      15'b000000000100000: n7949_o = n7941_o;
      15'b000000000010000: n7949_o = n7940_o;
      15'b000000000001000: n7949_o = n7939_o;
      15'b000000000000100: n7949_o = n7938_o;
      15'b000000000000010: n7949_o = n7937_o;
      15'b000000000000001: n7949_o = 4'b0000;
      default: n7949_o = 4'b0000;
    endcase
  /* control_mem_rtl.vhd:663:7  */
  assign n7951_o = s_bdata_mux == 4'b0000;
  assign n7952_o = psw[7];
  /* control_mem_rtl.vhd:664:44  */
  assign n7953_o = s_bit_data & n7952_o;
  /* control_mem_rtl.vhd:664:7  */
  assign n7955_o = s_bdata_mux == 4'b0001;
  /* control_mem_rtl.vhd:665:33  */
  assign n7956_o = ~s_bit_data;
  assign n7957_o = psw[7];
  /* control_mem_rtl.vhd:665:49  */
  assign n7958_o = n7956_o & n7957_o;
  /* control_mem_rtl.vhd:665:7  */
  assign n7960_o = s_bdata_mux == 4'b0010;
  /* control_mem_rtl.vhd:666:41  */
  assign n7961_o = new_cy_i[1];
  /* control_mem_rtl.vhd:666:7  */
  assign n7963_o = s_bdata_mux == 4'b0011;
  /* control_mem_rtl.vhd:667:7  */
  assign n7965_o = s_bdata_mux == 4'b0100;
  assign n7966_o = psw[7];
  /* control_mem_rtl.vhd:668:33  */
  assign n7967_o = ~n7966_o;
  /* control_mem_rtl.vhd:668:7  */
  assign n7969_o = s_bdata_mux == 4'b0101;
  /* control_mem_rtl.vhd:669:33  */
  assign n7970_o = ~s_bit_data;
  /* control_mem_rtl.vhd:669:7  */
  assign n7972_o = s_bdata_mux == 4'b0110;
  /* control_mem_rtl.vhd:670:7  */
  assign n7974_o = s_bdata_mux == 4'b0111;
  assign n7975_o = psw[7];
  /* control_mem_rtl.vhd:671:7  */
  assign n7977_o = s_bdata_mux == 4'b1000;
  assign n7978_o = psw[7];
  /* control_mem_rtl.vhd:672:44  */
  assign n7979_o = s_bit_data | n7978_o;
  /* control_mem_rtl.vhd:672:7  */
  assign n7981_o = s_bdata_mux == 4'b1001;
  /* control_mem_rtl.vhd:673:33  */
  assign n7982_o = ~s_bit_data;
  assign n7983_o = psw[7];
  /* control_mem_rtl.vhd:673:49  */
  assign n7984_o = n7982_o | n7983_o;
  /* control_mem_rtl.vhd:673:7  */
  assign n7986_o = s_bdata_mux == 4'b1010;
  /* control_mem_rtl.vhd:674:7  */
  assign n7988_o = s_bdata_mux == 4'b1011;
  assign n7989_o = {n7988_o, n7986_o, n7981_o, n7977_o, n7974_o, n7972_o, n7969_o, n7965_o, n7963_o, n7960_o, n7955_o, n7951_o};
  /* control_mem_rtl.vhd:662:5  */
  always @*
    case (n7989_o)
      12'b100000000000: n7993_o = 1'b1;
      12'b010000000000: n7993_o = n7984_o;
      12'b001000000000: n7993_o = n7979_o;
      12'b000100000000: n7993_o = n7975_o;
      12'b000010000000: n7993_o = s_bit_data;
      12'b000001000000: n7993_o = n7970_o;
      12'b000000100000: n7993_o = n7967_o;
      12'b000000010000: n7993_o = s_helpb;
      12'b000000001000: n7993_o = n7961_o;
      12'b000000000100: n7993_o = n7958_o;
      12'b000000000010: n7993_o = n7953_o;
      12'b000000000001: n7993_o = 1'b0;
      default: n7993_o = 1'b0;
    endcase
  /* control_mem_rtl.vhd:679:7  */
  assign n7995_o = s_adr_mux == 4'b0000;
  /* control_mem_rtl.vhd:680:7  */
  assign n7997_o = s_adr_mux == 4'b0001;
  /* control_mem_rtl.vhd:681:7  */
  assign n7999_o = s_adr_mux == 4'b0010;
  /* control_mem_rtl.vhd:682:7  */
  assign n8001_o = s_adr_mux == 4'b0011;
  /* control_mem_rtl.vhd:683:7  */
  assign n8003_o = s_adr_mux == 4'b0100;
  /* control_mem_rtl.vhd:684:7  */
  assign n8005_o = s_adr_mux == 4'b0101;
  /* control_mem_rtl.vhd:685:7  */
  assign n8007_o = s_adr_mux == 4'b0110;
  /* control_mem_rtl.vhd:686:7  */
  assign n8009_o = s_adr_mux == 4'b0111;
  /* control_mem_rtl.vhd:687:7  */
  assign n8011_o = s_adr_mux == 4'b1000;
  /* control_mem_rtl.vhd:688:7  */
  assign n8013_o = s_adr_mux == 4'b1001;
  /* control_mem_rtl.vhd:689:7  */
  assign n8015_o = s_adr_mux == 4'b1010;
  /* control_mem_rtl.vhd:690:7  */
  assign n8017_o = s_adr_mux == 4'b1011;
  /* control_mem_rtl.vhd:691:7  */
  assign n8019_o = s_adr_mux == 4'b1100;
  /* control_mem_rtl.vhd:692:7  */
  assign n8021_o = s_adr_mux == 4'b1101;
  /* control_mem_rtl.vhd:693:7  */
  assign n8023_o = s_adr_mux == 4'b1110;
  /* control_mem_rtl.vhd:694:34  */
  assign n8026_o = sp + 8'b00000001;
  /* control_mem_rtl.vhd:694:7  */
  assign n8028_o = s_adr_mux == 4'b1111;
  assign n8029_o = {n8028_o, n8023_o, n8021_o, n8019_o, n8017_o, n8015_o, n8013_o, n8011_o, n8009_o, n8007_o, n8005_o, n8003_o, n8001_o, n7999_o, n7997_o, n7995_o};
  /* control_mem_rtl.vhd:678:5  */
  always @*
    case (n8029_o)
      16'b1000000000000000: n8040_o = n8026_o;
      16'b0100000000000000: n8040_o = 8'b10000011;
      16'b0010000000000000: n8040_o = 8'b10000010;
      16'b0001000000000000: n8040_o = 8'b11110000;
      16'b0000100000000000: n8040_o = 8'b11010111;
      16'b0000010000000000: n8040_o = s_help;
      16'b0000001000000000: n8040_o = s_reg_data;
      16'b0000000100000000: n8040_o = rom_data_i;
      16'b0000000010000000: n8040_o = s_ri_data;
      16'b0000000001000000: n8040_o = s_rr_adr;
      16'b0000000000100000: n8040_o = sp;
      16'b0000000000010000: n8040_o = 8'b10001111;
      16'b0000000000001000: n8040_o = 8'b10001011;
      16'b0000000000000100: n8040_o = 8'b10001101;
      16'b0000000000000010: n8040_o = 8'b10001001;
      16'b0000000000000001: n8040_o = 8'b00000000;
      default: n8040_o = 8'b00000000;
    endcase
  /* control_mem_rtl.vhd:700:7  */
  assign n8042_o = s_adrx_mux == 2'b01;
  /* control_mem_rtl.vhd:704:7  */
  assign n8045_o = s_adrx_mux == 2'b10;
  assign n8046_o = {n8045_o, n8042_o};
  /* control_mem_rtl.vhd:698:5  */
  always @*
    case (n8046_o)
      2'b10: n8048_o = s_ri_data;
      2'b01: n8048_o = dpl;
      default: n8048_o = 8'b00000000;
    endcase
  /* control_mem_rtl.vhd:698:5  */
  always @*
    case (n8046_o)
      2'b10: n8050_o = 8'b00000000;
      2'b01: n8050_o = dph;
      default: n8050_o = 8'b00000000;
    endcase
  /* control_mem_rtl.vhd:698:5  */
  always @*
    case (n8046_o)
      2'b10: n8054_o = 1'b1;
      2'b01: n8054_o = 1'b1;
      default: n8054_o = 1'b0;
    endcase
  /* control_mem_rtl.vhd:712:7  */
  assign n8056_o = s_ri_adr == 8'b00000000;
  /* control_mem_rtl.vhd:713:7  */
  assign n8058_o = s_ri_adr == 8'b00000001;
  /* control_mem_rtl.vhd:714:7  */
  assign n8060_o = s_ri_adr == 8'b00001000;
  /* control_mem_rtl.vhd:715:7  */
  assign n8062_o = s_ri_adr == 8'b00001001;
  /* control_mem_rtl.vhd:716:7  */
  assign n8064_o = s_ri_adr == 8'b00010000;
  /* control_mem_rtl.vhd:717:7  */
  assign n8066_o = s_ri_adr == 8'b00010001;
  /* control_mem_rtl.vhd:718:7  */
  assign n8068_o = s_ri_adr == 8'b00011000;
  /* control_mem_rtl.vhd:719:7  */
  assign n8070_o = s_ri_adr == 8'b00011001;
  assign n8071_o = {n8070_o, n8068_o, n8066_o, n8064_o, n8062_o, n8060_o, n8058_o, n8056_o};
  /* control_mem_rtl.vhd:711:5  */
  always @*
    case (n8071_o)
      8'b10000000: n8073_o = s_r1_b3;
      8'b01000000: n8073_o = s_r0_b3;
      8'b00100000: n8073_o = s_r1_b2;
      8'b00010000: n8073_o = s_r0_b2;
      8'b00001000: n8073_o = s_r1_b1;
      8'b00000100: n8073_o = s_r0_b1;
      8'b00000010: n8073_o = s_r1_b0;
      8'b00000001: n8073_o = s_r0_b0;
      default: n8073_o = 8'b00000000;
    endcase
  /* control_mem_rtl.vhd:723:22  */
  assign n8075_o = s_regs_wr_en == 3'b100;
  /* control_mem_rtl.vhd:723:46  */
  assign n8077_o = s_regs_wr_en == 3'b101;
  /* control_mem_rtl.vhd:723:30  */
  assign n8078_o = n8075_o | n8077_o;
  /* control_mem_rtl.vhd:724:17  */
  assign n8079_o = s_adr[7];
  /* control_mem_rtl.vhd:725:37  */
  assign n8080_o = s_adr[7:4];
  /* control_mem_rtl.vhd:725:52  */
  assign n8082_o = n8080_o == 4'b0010;
  /* control_mem_rtl.vhd:724:26  */
  assign n8083_o = n8079_o | n8082_o;
  /* control_mem_rtl.vhd:726:38  */
  assign n8085_o = s_adr & 8'b11100110;
  /* control_mem_rtl.vhd:726:54  */
  assign n8087_o = n8085_o == 8'b00000000;
  /* control_mem_rtl.vhd:726:9  */
  assign n8088_o = n8083_o | n8087_o;
  /* control_mem_rtl.vhd:724:7  */
  assign n8091_o = n8088_o ? 1'b0 : 1'b1;
  /* control_mem_rtl.vhd:723:5  */
  assign n8093_o = n8078_o ? n8091_o : 1'b0;
  /* control_mem_rtl.vhd:772:17  */
  assign n8099_o = state == 3'b001;
  /* control_mem_rtl.vhd:777:11  */
  assign n8102_o = s_help_en == 4'b0000;
  /* control_mem_rtl.vhd:778:11  */
  assign n8104_o = s_help_en == 4'b0001;
  /* control_mem_rtl.vhd:779:11  */
  assign n8106_o = s_help_en == 4'b0010;
  /* control_mem_rtl.vhd:780:11  */
  assign n8108_o = s_help_en == 4'b0011;
  /* control_mem_rtl.vhd:781:11  */
  assign n8110_o = s_help_en == 4'b0100;
  /* control_mem_rtl.vhd:782:11  */
  assign n8112_o = s_help_en == 4'b0101;
  /* control_mem_rtl.vhd:783:11  */
  assign n8114_o = s_help_en == 4'b0110;
  /* control_mem_rtl.vhd:784:11  */
  assign n8116_o = s_help_en == 4'b0111;
  /* control_mem_rtl.vhd:785:11  */
  assign n8118_o = s_help_en == 4'b1000;
  /* control_mem_rtl.vhd:786:11  */
  assign n8120_o = s_help_en == 4'b1001;
  /* control_mem_rtl.vhd:787:11  */
  assign n8122_o = s_help_en == 4'b1010;
  assign n8123_o = {n8122_o, n8120_o, n8118_o, n8116_o, n8114_o, n8112_o, n8110_o, n8108_o, n8106_o, n8104_o, n8102_o};
  /* control_mem_rtl.vhd:776:9  */
  always @*
    case (n8123_o)
      11'b10000000000: n8129_o = acc;
      11'b01000000000: n8129_o = 8'b00100011;
      11'b00100000000: n8129_o = 8'b00011011;
      11'b00010000000: n8129_o = 8'b00010011;
      11'b00001000000: n8129_o = 8'b00001011;
      11'b00000100000: n8129_o = 8'b00000011;
      11'b00000010000: n8129_o = s_rr_adr;
      11'b00000001000: n8129_o = s_reg_data;
      11'b00000000100: n8129_o = aludata_i;
      11'b00000000010: n8129_o = rom_data_i;
      11'b00000000001: n8129_o = s_help;
      default: n8129_o = s_help;
    endcase
  /* control_mem_rtl.vhd:792:11  */
  assign n8131_o = s_help16_en == 2'b00;
  /* control_mem_rtl.vhd:793:39  */
  assign n8134_o = pc + 16'b0000000000000011;
  /* control_mem_rtl.vhd:793:11  */
  assign n8136_o = s_help16_en == 2'b01;
  /* control_mem_rtl.vhd:794:11  */
  assign n8138_o = s_help16_en == 2'b10;
  /* control_mem_rtl.vhd:795:11  */
  assign n8140_o = s_help16_en == 2'b11;
  assign n8141_o = {n8140_o, n8138_o, n8136_o, n8131_o};
  /* control_mem_rtl.vhd:791:9  */
  always @*
    case (n8141_o)
      4'b1000: n8142_o = pc_plus1;
      4'b0100: n8142_o = pc_plus2;
      4'b0010: n8142_o = n8134_o;
      4'b0001: n8142_o = s_help16;
      default: n8142_o = s_help16;
    endcase
  /* control_mem_rtl.vhd:800:11  */
  assign n8144_o = s_helpb_en == 1'b0;
  /* control_mem_rtl.vhd:801:42  */
  assign n8145_o = new_cy_i[1];
  /* control_mem_rtl.vhd:801:11  */
  assign n8147_o = s_helpb_en == 1'b1;
  assign n8148_o = {n8147_o, n8144_o};
  /* control_mem_rtl.vhd:799:9  */
  always @*
    case (n8148_o)
      2'b10: n8149_o = n8145_o;
      2'b01: n8149_o = s_helpb;
      default: n8149_o = s_helpb;
    endcase
  /* control_mem_rtl.vhd:863:7  */
  assign n8215_o = s_pc_inc_en == 4'b0001;
  /* control_mem_rtl.vhd:866:43  */
  assign n8216_o = {1'b0, pc_plus1};  //  uext
  /* control_mem_rtl.vhd:866:43  */
  assign n8217_o = {{9{rom_data_i[7]}}, rom_data_i}; // sext
  /* control_mem_rtl.vhd:866:43  */
  assign n8218_o = n8216_o + n8217_o;
  /* control_mem_rtl.vhd:866:20  */
  assign n8219_o = n8218_o[15:0];  // trunc
  /* control_mem_rtl.vhd:865:7  */
  assign n8221_o = s_pc_inc_en == 4'b0010;
  /* control_mem_rtl.vhd:867:7  */
  assign n8224_o = s_pc_inc_en == 4'b0011;
  /* control_mem_rtl.vhd:871:42  */
  assign n8225_o = s_help16[15:11];
  /* control_mem_rtl.vhd:872:37  */
  assign n8226_o = s_ir[7:5];
  /* control_mem_rtl.vhd:870:7  */
  assign n8228_o = s_pc_inc_en == 4'b0100;
  assign n8229_o = {dph, dpl};
  /* control_mem_rtl.vhd:875:27  */
  assign n8230_o = {8'b0, acc};  //  uext
  /* control_mem_rtl.vhd:875:27  */
  assign n8231_o = n8229_o + n8230_o;
  /* control_mem_rtl.vhd:874:7  */
  assign n8233_o = s_pc_inc_en == 4'b0101;
  /* control_mem_rtl.vhd:876:7  */
  assign n8235_o = s_pc_inc_en == 4'b0110;
  /* control_mem_rtl.vhd:878:7  */
  assign n8237_o = s_pc_inc_en == 4'b0111;
  /* control_mem_rtl.vhd:881:7  */
  assign n8239_o = s_pc_inc_en == 4'b1000;
  /* control_mem_rtl.vhd:885:29  */
  assign n8240_o = {8'b0, acc};  //  uext
  /* control_mem_rtl.vhd:885:29  */
  assign n8241_o = pc_plus1 + n8240_o;
  /* control_mem_rtl.vhd:884:7  */
  assign n8243_o = s_pc_inc_en == 4'b1001;
  assign n8244_o = {n8243_o, n8239_o, n8237_o, n8235_o, n8233_o, n8228_o, n8224_o, n8221_o, n8215_o};
  assign n8245_o = pc_plus1[7:0];
  assign n8246_o = n8219_o[7:0];
  assign n8247_o = n8231_o[7:0];
  assign n8248_o = s_help16[7:0];
  assign n8249_o = n8241_o[7:0];
  assign n8250_o = pc[7:0];
  /* control_mem_rtl.vhd:862:5  */
  always @*
    case (n8244_o)
      9'b100000000: n8251_o = n8249_o;
      9'b010000000: n8251_o = s_reg_data;
      9'b001000000: n8251_o = rom_data_i;
      9'b000100000: n8251_o = n8248_o;
      9'b000010000: n8251_o = n8247_o;
      9'b000001000: n8251_o = rom_data_i;
      9'b000000100: n8251_o = s_help;
      9'b000000010: n8251_o = n8246_o;
      9'b000000001: n8251_o = n8245_o;
      default: n8251_o = n8250_o;
    endcase
  assign n8252_o = pc_plus1[10:8];
  assign n8253_o = n8219_o[10:8];
  assign n8254_o = n8222_o[2:0];
  assign n8255_o = n8231_o[10:8];
  assign n8256_o = s_help16[10:8];
  assign n8257_o = s_help[2:0];
  assign n8258_o = s_help[2:0];
  assign n8259_o = n8241_o[10:8];
  assign n8260_o = pc[10:8];
  /* control_mem_rtl.vhd:862:5  */
  always @*
    case (n8244_o)
      9'b100000000: n8261_o = n8259_o;
      9'b010000000: n8261_o = n8258_o;
      9'b001000000: n8261_o = n8257_o;
      9'b000100000: n8261_o = n8256_o;
      9'b000010000: n8261_o = n8255_o;
      9'b000001000: n8261_o = n8226_o;
      9'b000000100: n8261_o = n8254_o;
      9'b000000010: n8261_o = n8253_o;
      9'b000000001: n8261_o = n8252_o;
      default: n8261_o = n8260_o;
    endcase
  assign n8262_o = pc_plus1[15:11];
  assign n8263_o = n8219_o[15:11];
  assign n8264_o = n8222_o[7:3];
  assign n8265_o = n8231_o[15:11];
  assign n8266_o = s_help16[15:11];
  assign n8267_o = s_help[7:3];
  assign n8268_o = s_help[7:3];
  assign n8269_o = n8241_o[15:11];
  assign n8270_o = pc[15:11];
  /* control_mem_rtl.vhd:862:5  */
  always @*
    case (n8244_o)
      9'b100000000: n8271_o = n8269_o;
      9'b010000000: n8271_o = n8268_o;
      9'b001000000: n8271_o = n8267_o;
      9'b000100000: n8271_o = n8266_o;
      9'b000010000: n8271_o = n8265_o;
      9'b000001000: n8271_o = n8225_o;
      9'b000000100: n8271_o = n8264_o;
      9'b000000010: n8271_o = n8263_o;
      9'b000000001: n8271_o = n8262_o;
      default: n8271_o = n8270_o;
    endcase
  /* control_mem_rtl.vhd:956:32  */
  assign n8293_o = tcon[3];
  /* control_mem_rtl.vhd:956:48  */
  assign n8294_o = tcon[2];
  /* control_mem_rtl.vhd:956:52  */
  assign n8295_o = n8294_o & s_int1_edge;
  /* control_mem_rtl.vhd:957:38  */
  assign n8296_o = tcon[2];
  /* control_mem_rtl.vhd:957:27  */
  assign n8297_o = ~n8296_o;
  /* control_mem_rtl.vhd:957:46  */
  assign n8298_o = ~s_int1_h2;
  /* control_mem_rtl.vhd:957:42  */
  assign n8299_o = n8297_o & n8298_o;
  /* control_mem_rtl.vhd:958:42  */
  assign n8300_o = s_ext1isr_d | s_ext1isrh_d;
  /* control_mem_rtl.vhd:958:26  */
  assign n8301_o = ~n8300_o;
  /* control_mem_rtl.vhd:957:64  */
  assign n8302_o = n8299_o & n8301_o;
  /* control_mem_rtl.vhd:956:72  */
  assign n8303_o = n8295_o | n8302_o;
  /* control_mem_rtl.vhd:956:36  */
  assign n8304_o = n8293_o | n8303_o;
  /* control_mem_rtl.vhd:959:32  */
  assign n8305_o = tcon[1];
  /* control_mem_rtl.vhd:959:48  */
  assign n8306_o = tcon[0];
  /* control_mem_rtl.vhd:959:52  */
  assign n8307_o = n8306_o & s_int0_edge;
  /* control_mem_rtl.vhd:960:38  */
  assign n8308_o = tcon[0];
  /* control_mem_rtl.vhd:960:27  */
  assign n8309_o = ~n8308_o;
  /* control_mem_rtl.vhd:960:46  */
  assign n8310_o = ~s_int0_h2;
  /* control_mem_rtl.vhd:960:42  */
  assign n8311_o = n8309_o & n8310_o;
  /* control_mem_rtl.vhd:961:42  */
  assign n8312_o = s_ext0isr_d | s_ext0isrh_d;
  /* control_mem_rtl.vhd:961:26  */
  assign n8313_o = ~n8312_o;
  /* control_mem_rtl.vhd:960:64  */
  assign n8314_o = n8311_o & n8313_o;
  /* control_mem_rtl.vhd:959:72  */
  assign n8315_o = n8307_o | n8314_o;
  /* control_mem_rtl.vhd:959:36  */
  assign n8316_o = n8305_o | n8315_o;
  /* control_mem_rtl.vhd:962:32  */
  assign n8317_o = tcon[5];
  /* control_mem_rtl.vhd:962:36  */
  assign n8318_o = n8317_o | s_tf0_edge;
  /* control_mem_rtl.vhd:963:32  */
  assign n8319_o = tcon[7];
  /* control_mem_rtl.vhd:963:36  */
  assign n8320_o = n8319_o | s_tf1_edge;
  /* control_mem_rtl.vhd:967:32  */
  assign n8321_o = scon[0];
  /* control_mem_rtl.vhd:967:36  */
  assign n8322_o = n8321_o | s_ri_edge;
  /* control_mem_rtl.vhd:968:32  */
  assign n8323_o = scon[1];
  /* control_mem_rtl.vhd:968:36  */
  assign n8324_o = n8323_o | s_ti_edge;
  /* control_mem_rtl.vhd:974:27  */
  assign n8325_o = ~s_intblock;
  /* control_mem_rtl.vhd:974:32  */
  assign n8326_o = n8325_o & s_intpre;
  /* control_mem_rtl.vhd:974:58  */
  assign n8328_o = state == 3'b001;
  /* control_mem_rtl.vhd:974:49  */
  assign n8329_o = n8326_o & n8328_o;
  /* control_mem_rtl.vhd:974:66  */
  assign n8330_o = n8329_o | s_intpre2;
  /* control_mem_rtl.vhd:975:24  */
  assign n8333_o = sp + 8'b00000001;
  /* control_mem_rtl.vhd:979:28  */
  assign n8336_o = sp - 8'b00000001;
  /* control_mem_rtl.vhd:978:17  */
  assign n8338_o = s_command == 8'b00100010;
  /* control_mem_rtl.vhd:978:26  */
  assign n8340_o = s_command == 8'b00110010;
  /* control_mem_rtl.vhd:978:26  */
  assign n8341_o = n8338_o | n8340_o;
  /* control_mem_rtl.vhd:981:28  */
  assign n8344_o = sp + 8'b00000001;
  /* control_mem_rtl.vhd:977:15  */
  always @*
    case (n8341_o)
      1'b1: n8345_o = n8336_o;
      default: n8345_o = n8344_o;
    endcase
  /* control_mem_rtl.vhd:974:13  */
  assign n8346_o = n8330_o ? n8333_o : n8345_o;
  /* control_mem_rtl.vhd:972:11  */
  assign n8348_o = s_regs_wr_en == 3'b001;
  /* control_mem_rtl.vhd:984:11  */
  assign n8350_o = s_regs_wr_en == 3'b010;
  /* control_mem_rtl.vhd:988:31  */
  assign n8351_o = new_cy_i[1];
  /* control_mem_rtl.vhd:989:31  */
  assign n8352_o = new_cy_i[0];
  /* control_mem_rtl.vhd:986:11  */
  assign n8354_o = s_regs_wr_en == 3'b011;
  /* control_mem_rtl.vhd:994:20  */
  assign n8355_o = {24'b0, s_adr};  //  uext
  /* control_mem_rtl.vhd:994:40  */
  assign n8357_o = n8355_o == 32'b00000000000000000000000010000001;
  /* control_mem_rtl.vhd:994:17  */
  assign n8358_o = n8357_o ? s_data : sp;
  /* control_mem_rtl.vhd:993:15  */
  assign n8360_o = s_regs_wr_en == 3'b100;
  /* control_mem_rtl.vhd:998:31  */
  assign n8361_o = ~s_intblock;
  /* control_mem_rtl.vhd:998:36  */
  assign n8362_o = n8361_o & s_intpre;
  /* control_mem_rtl.vhd:998:62  */
  assign n8364_o = state == 3'b001;
  /* control_mem_rtl.vhd:998:53  */
  assign n8365_o = n8362_o & n8364_o;
  /* control_mem_rtl.vhd:998:70  */
  assign n8366_o = n8365_o | s_intpre2;
  /* control_mem_rtl.vhd:999:28  */
  assign n8369_o = sp + 8'b00000001;
  /* control_mem_rtl.vhd:1001:32  */
  assign n8371_o = s_command == 8'b11010000;
  /* control_mem_rtl.vhd:1002:25  */
  assign n8372_o = {24'b0, s_adr};  //  uext
  /* control_mem_rtl.vhd:1002:45  */
  assign n8374_o = n8372_o == 32'b00000000000000000000000010000001;
  /* control_mem_rtl.vhd:1005:32  */
  assign n8377_o = sp - 8'b00000001;
  /* control_mem_rtl.vhd:1002:21  */
  assign n8378_o = n8374_o ? s_data : n8377_o;
  /* control_mem_rtl.vhd:1008:30  */
  assign n8381_o = sp + 8'b00000001;
  /* control_mem_rtl.vhd:1001:19  */
  assign n8382_o = n8371_o ? n8378_o : n8381_o;
  /* control_mem_rtl.vhd:998:17  */
  assign n8383_o = n8366_o ? n8369_o : n8382_o;
  /* control_mem_rtl.vhd:997:15  */
  assign n8385_o = s_regs_wr_en == 3'b101;
  assign n8386_o = {n8385_o, n8360_o};
  /* control_mem_rtl.vhd:992:13  */
  always @*
    case (n8386_o)
      2'b10: n8387_o = n8383_o;
      2'b01: n8387_o = n8358_o;
      default: n8387_o = sp;
    endcase
  /* control_mem_rtl.vhd:1014:21  */
  assign n8388_o = s_adr[7];
  /* control_mem_rtl.vhd:1015:20  */
  assign n8389_o = {24'b0, s_adr};  //  uext
  /* control_mem_rtl.vhd:1016:15  */
  assign n8391_o = n8389_o == 32'b00000000000000000000000010000000;
  /* control_mem_rtl.vhd:1017:15  */
  assign n8393_o = n8389_o == 32'b00000000000000000000000010000010;
  /* control_mem_rtl.vhd:1018:15  */
  assign n8395_o = n8389_o == 32'b00000000000000000000000010000011;
  /* control_mem_rtl.vhd:1020:31  */
  assign n8396_o = s_data[3:0];
  /* control_mem_rtl.vhd:1021:44  */
  assign n8397_o = s_data[7];
  /* control_mem_rtl.vhd:1019:15  */
  assign n8399_o = n8389_o == 32'b00000000000000000000000010000111;
  /* control_mem_rtl.vhd:1022:15  */
  assign n8401_o = n8389_o == 32'b00000000000000000000000010001000;
  /* control_mem_rtl.vhd:1023:15  */
  assign n8403_o = n8389_o == 32'b00000000000000000000000010001001;
  /* control_mem_rtl.vhd:1024:15  */
  assign n8405_o = n8389_o == 32'b00000000000000000000000010001010;
  /* control_mem_rtl.vhd:1028:15  */
  assign n8407_o = n8389_o == 32'b00000000000000000000000010001011;
  /* control_mem_rtl.vhd:1032:15  */
  assign n8409_o = n8389_o == 32'b00000000000000000000000010001100;
  /* control_mem_rtl.vhd:1036:15  */
  assign n8411_o = n8389_o == 32'b00000000000000000000000010001101;
  /* control_mem_rtl.vhd:1040:15  */
  assign n8413_o = n8389_o == 32'b00000000000000000000000010001110;
  /* control_mem_rtl.vhd:1041:15  */
  assign n8415_o = n8389_o == 32'b00000000000000000000000010010000;
  /* control_mem_rtl.vhd:1042:15  */
  assign n8417_o = n8389_o == 32'b00000000000000000000000010011000;
  /* control_mem_rtl.vhd:1043:15  */
  assign n8419_o = n8389_o == 32'b00000000000000000000000010011001;
  /* control_mem_rtl.vhd:1046:15  */
  assign n8421_o = n8389_o == 32'b00000000000000000000000010011010;
  /* control_mem_rtl.vhd:1047:15  */
  assign n8423_o = n8389_o == 32'b00000000000000000000000010100000;
  /* control_mem_rtl.vhd:1048:15  */
  assign n8425_o = n8389_o == 32'b00000000000000000000000010101000;
  /* control_mem_rtl.vhd:1049:15  */
  assign n8427_o = n8389_o == 32'b00000000000000000000000010110000;
  /* control_mem_rtl.vhd:1050:15  */
  assign n8429_o = n8389_o == 32'b00000000000000000000000010111000;
  /* control_mem_rtl.vhd:1052:64  */
  assign n8430_o = s_data[7:1];
  /* control_mem_rtl.vhd:1051:15  */
  assign n8432_o = n8389_o == 32'b00000000000000000000000011010000;
  /* control_mem_rtl.vhd:1053:15  */
  assign n8434_o = n8389_o == 32'b00000000000000000000000011100000;
  /* control_mem_rtl.vhd:1054:15  */
  assign n8436_o = n8389_o == 32'b00000000000000000000000011110000;
  assign n8437_o = {n8436_o, n8434_o, n8432_o, n8429_o, n8427_o, n8425_o, n8423_o, n8421_o, n8419_o, n8417_o, n8415_o, n8413_o, n8411_o, n8409_o, n8407_o, n8405_o, n8403_o, n8401_o, n8399_o, n8395_o, n8393_o, n8391_o};
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8440_o = 1'b0;
      22'b0100000000000000000000: n8440_o = 1'b0;
      22'b0010000000000000000000: n8440_o = 1'b0;
      22'b0001000000000000000000: n8440_o = 1'b0;
      22'b0000100000000000000000: n8440_o = 1'b0;
      22'b0000010000000000000000: n8440_o = 1'b0;
      22'b0000001000000000000000: n8440_o = 1'b0;
      22'b0000000100000000000000: n8440_o = 1'b0;
      22'b0000000010000000000000: n8440_o = 1'b1;
      22'b0000000001000000000000: n8440_o = 1'b0;
      22'b0000000000100000000000: n8440_o = 1'b0;
      22'b0000000000010000000000: n8440_o = 1'b0;
      22'b0000000000001000000000: n8440_o = 1'b0;
      22'b0000000000000100000000: n8440_o = 1'b0;
      22'b0000000000000010000000: n8440_o = 1'b0;
      22'b0000000000000001000000: n8440_o = 1'b0;
      22'b0000000000000000100000: n8440_o = 1'b0;
      22'b0000000000000000010000: n8440_o = 1'b0;
      22'b0000000000000000001000: n8440_o = 1'b0;
      22'b0000000000000000000100: n8440_o = 1'b0;
      22'b0000000000000000000010: n8440_o = 1'b0;
      22'b0000000000000000000001: n8440_o = 1'b0;
      default: n8440_o = 1'b0;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8446_o = 1'b0;
      22'b0100000000000000000000: n8446_o = 1'b0;
      22'b0010000000000000000000: n8446_o = 1'b0;
      22'b0001000000000000000000: n8446_o = 1'b0;
      22'b0000100000000000000000: n8446_o = 1'b0;
      22'b0000010000000000000000: n8446_o = 1'b0;
      22'b0000001000000000000000: n8446_o = 1'b0;
      22'b0000000100000000000000: n8446_o = 1'b0;
      22'b0000000010000000000000: n8446_o = 1'b0;
      22'b0000000001000000000000: n8446_o = 1'b0;
      22'b0000000000100000000000: n8446_o = 1'b0;
      22'b0000000000010000000000: n8446_o = 1'b0;
      22'b0000000000001000000000: n8446_o = 1'b1;
      22'b0000000000000100000000: n8446_o = 1'b1;
      22'b0000000000000010000000: n8446_o = 1'b1;
      22'b0000000000000001000000: n8446_o = 1'b1;
      22'b0000000000000000100000: n8446_o = 1'b0;
      22'b0000000000000000010000: n8446_o = 1'b0;
      22'b0000000000000000001000: n8446_o = 1'b0;
      22'b0000000000000000000100: n8446_o = 1'b0;
      22'b0000000000000000000010: n8446_o = 1'b0;
      22'b0000000000000000000001: n8446_o = 1'b0;
      default: n8446_o = 1'b0;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8447_o = s_smodreg;
      22'b0100000000000000000000: n8447_o = s_smodreg;
      22'b0010000000000000000000: n8447_o = s_smodreg;
      22'b0001000000000000000000: n8447_o = s_smodreg;
      22'b0000100000000000000000: n8447_o = s_smodreg;
      22'b0000010000000000000000: n8447_o = s_smodreg;
      22'b0000001000000000000000: n8447_o = s_smodreg;
      22'b0000000100000000000000: n8447_o = s_smodreg;
      22'b0000000010000000000000: n8447_o = s_smodreg;
      22'b0000000001000000000000: n8447_o = s_smodreg;
      22'b0000000000100000000000: n8447_o = s_smodreg;
      22'b0000000000010000000000: n8447_o = s_smodreg;
      22'b0000000000001000000000: n8447_o = s_smodreg;
      22'b0000000000000100000000: n8447_o = s_smodreg;
      22'b0000000000000010000000: n8447_o = s_smodreg;
      22'b0000000000000001000000: n8447_o = s_smodreg;
      22'b0000000000000000100000: n8447_o = s_smodreg;
      22'b0000000000000000010000: n8447_o = s_smodreg;
      22'b0000000000000000001000: n8447_o = n8397_o;
      22'b0000000000000000000100: n8447_o = s_smodreg;
      22'b0000000000000000000010: n8447_o = s_smodreg;
      22'b0000000000000000000001: n8447_o = s_smodreg;
      default: n8447_o = s_smodreg;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8448_o = s_reload;
      22'b0100000000000000000000: n8448_o = s_reload;
      22'b0010000000000000000000: n8448_o = s_reload;
      22'b0001000000000000000000: n8448_o = s_reload;
      22'b0000100000000000000000: n8448_o = s_reload;
      22'b0000010000000000000000: n8448_o = s_reload;
      22'b0000001000000000000000: n8448_o = s_reload;
      22'b0000000100000000000000: n8448_o = s_reload;
      22'b0000000010000000000000: n8448_o = s_reload;
      22'b0000000001000000000000: n8448_o = s_reload;
      22'b0000000000100000000000: n8448_o = s_reload;
      22'b0000000000010000000000: n8448_o = s_reload;
      22'b0000000000001000000000: n8448_o = s_data;
      22'b0000000000000100000000: n8448_o = s_data;
      22'b0000000000000010000000: n8448_o = s_data;
      22'b0000000000000001000000: n8448_o = s_data;
      22'b0000000000000000100000: n8448_o = s_reload;
      22'b0000000000000000010000: n8448_o = s_reload;
      22'b0000000000000000001000: n8448_o = s_reload;
      22'b0000000000000000000100: n8448_o = s_reload;
      22'b0000000000000000000010: n8448_o = s_reload;
      22'b0000000000000000000001: n8448_o = s_reload;
      default: n8448_o = s_reload;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8453_o = s_wt;
      22'b0100000000000000000000: n8453_o = s_wt;
      22'b0010000000000000000000: n8453_o = s_wt;
      22'b0001000000000000000000: n8453_o = s_wt;
      22'b0000100000000000000000: n8453_o = s_wt;
      22'b0000010000000000000000: n8453_o = s_wt;
      22'b0000001000000000000000: n8453_o = s_wt;
      22'b0000000100000000000000: n8453_o = s_wt;
      22'b0000000010000000000000: n8453_o = s_wt;
      22'b0000000001000000000000: n8453_o = s_wt;
      22'b0000000000100000000000: n8453_o = s_wt;
      22'b0000000000010000000000: n8453_o = s_wt;
      22'b0000000000001000000000: n8453_o = 2'b11;
      22'b0000000000000100000000: n8453_o = 2'b10;
      22'b0000000000000010000000: n8453_o = 2'b01;
      22'b0000000000000001000000: n8453_o = 2'b00;
      22'b0000000000000000100000: n8453_o = s_wt;
      22'b0000000000000000010000: n8453_o = s_wt;
      22'b0000000000000000001000: n8453_o = s_wt;
      22'b0000000000000000000100: n8453_o = s_wt;
      22'b0000000000000000000010: n8453_o = s_wt;
      22'b0000000000000000000001: n8453_o = s_wt;
      default: n8453_o = s_wt;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8454_o = p0;
      22'b0100000000000000000000: n8454_o = p0;
      22'b0010000000000000000000: n8454_o = p0;
      22'b0001000000000000000000: n8454_o = p0;
      22'b0000100000000000000000: n8454_o = p0;
      22'b0000010000000000000000: n8454_o = p0;
      22'b0000001000000000000000: n8454_o = p0;
      22'b0000000100000000000000: n8454_o = p0;
      22'b0000000010000000000000: n8454_o = p0;
      22'b0000000001000000000000: n8454_o = p0;
      22'b0000000000100000000000: n8454_o = p0;
      22'b0000000000010000000000: n8454_o = p0;
      22'b0000000000001000000000: n8454_o = p0;
      22'b0000000000000100000000: n8454_o = p0;
      22'b0000000000000010000000: n8454_o = p0;
      22'b0000000000000001000000: n8454_o = p0;
      22'b0000000000000000100000: n8454_o = p0;
      22'b0000000000000000010000: n8454_o = p0;
      22'b0000000000000000001000: n8454_o = p0;
      22'b0000000000000000000100: n8454_o = p0;
      22'b0000000000000000000010: n8454_o = p0;
      22'b0000000000000000000001: n8454_o = s_data;
      default: n8454_o = p0;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8455_o = dpl;
      22'b0100000000000000000000: n8455_o = dpl;
      22'b0010000000000000000000: n8455_o = dpl;
      22'b0001000000000000000000: n8455_o = dpl;
      22'b0000100000000000000000: n8455_o = dpl;
      22'b0000010000000000000000: n8455_o = dpl;
      22'b0000001000000000000000: n8455_o = dpl;
      22'b0000000100000000000000: n8455_o = dpl;
      22'b0000000010000000000000: n8455_o = dpl;
      22'b0000000001000000000000: n8455_o = dpl;
      22'b0000000000100000000000: n8455_o = dpl;
      22'b0000000000010000000000: n8455_o = dpl;
      22'b0000000000001000000000: n8455_o = dpl;
      22'b0000000000000100000000: n8455_o = dpl;
      22'b0000000000000010000000: n8455_o = dpl;
      22'b0000000000000001000000: n8455_o = dpl;
      22'b0000000000000000100000: n8455_o = dpl;
      22'b0000000000000000010000: n8455_o = dpl;
      22'b0000000000000000001000: n8455_o = dpl;
      22'b0000000000000000000100: n8455_o = dpl;
      22'b0000000000000000000010: n8455_o = s_data;
      22'b0000000000000000000001: n8455_o = dpl;
      default: n8455_o = dpl;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8456_o = dph;
      22'b0100000000000000000000: n8456_o = dph;
      22'b0010000000000000000000: n8456_o = dph;
      22'b0001000000000000000000: n8456_o = dph;
      22'b0000100000000000000000: n8456_o = dph;
      22'b0000010000000000000000: n8456_o = dph;
      22'b0000001000000000000000: n8456_o = dph;
      22'b0000000100000000000000: n8456_o = dph;
      22'b0000000010000000000000: n8456_o = dph;
      22'b0000000001000000000000: n8456_o = dph;
      22'b0000000000100000000000: n8456_o = dph;
      22'b0000000000010000000000: n8456_o = dph;
      22'b0000000000001000000000: n8456_o = dph;
      22'b0000000000000100000000: n8456_o = dph;
      22'b0000000000000010000000: n8456_o = dph;
      22'b0000000000000001000000: n8456_o = dph;
      22'b0000000000000000100000: n8456_o = dph;
      22'b0000000000000000010000: n8456_o = dph;
      22'b0000000000000000001000: n8456_o = dph;
      22'b0000000000000000000100: n8456_o = s_data;
      22'b0000000000000000000010: n8456_o = dph;
      22'b0000000000000000000001: n8456_o = dph;
      default: n8456_o = dph;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8457_o = pcon;
      22'b0100000000000000000000: n8457_o = pcon;
      22'b0010000000000000000000: n8457_o = pcon;
      22'b0001000000000000000000: n8457_o = pcon;
      22'b0000100000000000000000: n8457_o = pcon;
      22'b0000010000000000000000: n8457_o = pcon;
      22'b0000001000000000000000: n8457_o = pcon;
      22'b0000000100000000000000: n8457_o = pcon;
      22'b0000000010000000000000: n8457_o = pcon;
      22'b0000000001000000000000: n8457_o = pcon;
      22'b0000000000100000000000: n8457_o = pcon;
      22'b0000000000010000000000: n8457_o = pcon;
      22'b0000000000001000000000: n8457_o = pcon;
      22'b0000000000000100000000: n8457_o = pcon;
      22'b0000000000000010000000: n8457_o = pcon;
      22'b0000000000000001000000: n8457_o = pcon;
      22'b0000000000000000100000: n8457_o = pcon;
      22'b0000000000000000010000: n8457_o = pcon;
      22'b0000000000000000001000: n8457_o = n8396_o;
      22'b0000000000000000000100: n8457_o = pcon;
      22'b0000000000000000000010: n8457_o = pcon;
      22'b0000000000000000000001: n8457_o = pcon;
      default: n8457_o = pcon;
    endcase
  assign n8458_o = tcon[0];
  assign n8459_o = tcon[2];
  assign n8460_o = tcon[4];
  assign n8461_o = tcon[6];
  assign n8462_o = {n8320_o, n8461_o, n8318_o, n8460_o, n8304_o, n8459_o, n8316_o, n8458_o};
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8463_o = n8462_o;
      22'b0100000000000000000000: n8463_o = n8462_o;
      22'b0010000000000000000000: n8463_o = n8462_o;
      22'b0001000000000000000000: n8463_o = n8462_o;
      22'b0000100000000000000000: n8463_o = n8462_o;
      22'b0000010000000000000000: n8463_o = n8462_o;
      22'b0000001000000000000000: n8463_o = n8462_o;
      22'b0000000100000000000000: n8463_o = n8462_o;
      22'b0000000010000000000000: n8463_o = n8462_o;
      22'b0000000001000000000000: n8463_o = n8462_o;
      22'b0000000000100000000000: n8463_o = n8462_o;
      22'b0000000000010000000000: n8463_o = n8462_o;
      22'b0000000000001000000000: n8463_o = n8462_o;
      22'b0000000000000100000000: n8463_o = n8462_o;
      22'b0000000000000010000000: n8463_o = n8462_o;
      22'b0000000000000001000000: n8463_o = n8462_o;
      22'b0000000000000000100000: n8463_o = n8462_o;
      22'b0000000000000000010000: n8463_o = s_data;
      22'b0000000000000000001000: n8463_o = n8462_o;
      22'b0000000000000000000100: n8463_o = n8462_o;
      22'b0000000000000000000010: n8463_o = n8462_o;
      22'b0000000000000000000001: n8463_o = n8462_o;
      default: n8463_o = n8462_o;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8464_o = tmod;
      22'b0100000000000000000000: n8464_o = tmod;
      22'b0010000000000000000000: n8464_o = tmod;
      22'b0001000000000000000000: n8464_o = tmod;
      22'b0000100000000000000000: n8464_o = tmod;
      22'b0000010000000000000000: n8464_o = tmod;
      22'b0000001000000000000000: n8464_o = tmod;
      22'b0000000100000000000000: n8464_o = tmod;
      22'b0000000010000000000000: n8464_o = tmod;
      22'b0000000001000000000000: n8464_o = tmod;
      22'b0000000000100000000000: n8464_o = tmod;
      22'b0000000000010000000000: n8464_o = tmod;
      22'b0000000000001000000000: n8464_o = tmod;
      22'b0000000000000100000000: n8464_o = tmod;
      22'b0000000000000010000000: n8464_o = tmod;
      22'b0000000000000001000000: n8464_o = tmod;
      22'b0000000000000000100000: n8464_o = s_data;
      22'b0000000000000000010000: n8464_o = tmod;
      22'b0000000000000000001000: n8464_o = tmod;
      22'b0000000000000000000100: n8464_o = tmod;
      22'b0000000000000000000010: n8464_o = tmod;
      22'b0000000000000000000001: n8464_o = tmod;
      default: n8464_o = tmod;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8465_o = p1;
      22'b0100000000000000000000: n8465_o = p1;
      22'b0010000000000000000000: n8465_o = p1;
      22'b0001000000000000000000: n8465_o = p1;
      22'b0000100000000000000000: n8465_o = p1;
      22'b0000010000000000000000: n8465_o = p1;
      22'b0000001000000000000000: n8465_o = p1;
      22'b0000000100000000000000: n8465_o = p1;
      22'b0000000010000000000000: n8465_o = p1;
      22'b0000000001000000000000: n8465_o = p1;
      22'b0000000000100000000000: n8465_o = s_data;
      22'b0000000000010000000000: n8465_o = p1;
      22'b0000000000001000000000: n8465_o = p1;
      22'b0000000000000100000000: n8465_o = p1;
      22'b0000000000000010000000: n8465_o = p1;
      22'b0000000000000001000000: n8465_o = p1;
      22'b0000000000000000100000: n8465_o = p1;
      22'b0000000000000000010000: n8465_o = p1;
      22'b0000000000000000001000: n8465_o = p1;
      22'b0000000000000000000100: n8465_o = p1;
      22'b0000000000000000000010: n8465_o = p1;
      22'b0000000000000000000001: n8465_o = p1;
      default: n8465_o = p1;
    endcase
  assign n8466_o = scon[7:2];
  assign n8467_o = {n8466_o, n8324_o, n8322_o};
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8468_o = n8467_o;
      22'b0100000000000000000000: n8468_o = n8467_o;
      22'b0010000000000000000000: n8468_o = n8467_o;
      22'b0001000000000000000000: n8468_o = n8467_o;
      22'b0000100000000000000000: n8468_o = n8467_o;
      22'b0000010000000000000000: n8468_o = n8467_o;
      22'b0000001000000000000000: n8468_o = n8467_o;
      22'b0000000100000000000000: n8468_o = n8467_o;
      22'b0000000010000000000000: n8468_o = n8467_o;
      22'b0000000001000000000000: n8468_o = s_data;
      22'b0000000000100000000000: n8468_o = n8467_o;
      22'b0000000000010000000000: n8468_o = n8467_o;
      22'b0000000000001000000000: n8468_o = n8467_o;
      22'b0000000000000100000000: n8468_o = n8467_o;
      22'b0000000000000010000000: n8468_o = n8467_o;
      22'b0000000000000001000000: n8468_o = n8467_o;
      22'b0000000000000000100000: n8468_o = n8467_o;
      22'b0000000000000000010000: n8468_o = n8467_o;
      22'b0000000000000000001000: n8468_o = n8467_o;
      22'b0000000000000000000100: n8468_o = n8467_o;
      22'b0000000000000000000010: n8468_o = n8467_o;
      22'b0000000000000000000001: n8468_o = n8467_o;
      default: n8468_o = n8467_o;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8469_o = sbuf;
      22'b0100000000000000000000: n8469_o = sbuf;
      22'b0010000000000000000000: n8469_o = sbuf;
      22'b0001000000000000000000: n8469_o = sbuf;
      22'b0000100000000000000000: n8469_o = sbuf;
      22'b0000010000000000000000: n8469_o = sbuf;
      22'b0000001000000000000000: n8469_o = sbuf;
      22'b0000000100000000000000: n8469_o = sbuf;
      22'b0000000010000000000000: n8469_o = s_data;
      22'b0000000001000000000000: n8469_o = sbuf;
      22'b0000000000100000000000: n8469_o = sbuf;
      22'b0000000000010000000000: n8469_o = sbuf;
      22'b0000000000001000000000: n8469_o = sbuf;
      22'b0000000000000100000000: n8469_o = sbuf;
      22'b0000000000000010000000: n8469_o = sbuf;
      22'b0000000000000001000000: n8469_o = sbuf;
      22'b0000000000000000100000: n8469_o = sbuf;
      22'b0000000000000000010000: n8469_o = sbuf;
      22'b0000000000000000001000: n8469_o = sbuf;
      22'b0000000000000000000100: n8469_o = sbuf;
      22'b0000000000000000000010: n8469_o = sbuf;
      22'b0000000000000000000001: n8469_o = sbuf;
      default: n8469_o = sbuf;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8470_o = p2;
      22'b0100000000000000000000: n8470_o = p2;
      22'b0010000000000000000000: n8470_o = p2;
      22'b0001000000000000000000: n8470_o = p2;
      22'b0000100000000000000000: n8470_o = p2;
      22'b0000010000000000000000: n8470_o = p2;
      22'b0000001000000000000000: n8470_o = s_data;
      22'b0000000100000000000000: n8470_o = p2;
      22'b0000000010000000000000: n8470_o = p2;
      22'b0000000001000000000000: n8470_o = p2;
      22'b0000000000100000000000: n8470_o = p2;
      22'b0000000000010000000000: n8470_o = p2;
      22'b0000000000001000000000: n8470_o = p2;
      22'b0000000000000100000000: n8470_o = p2;
      22'b0000000000000010000000: n8470_o = p2;
      22'b0000000000000001000000: n8470_o = p2;
      22'b0000000000000000100000: n8470_o = p2;
      22'b0000000000000000010000: n8470_o = p2;
      22'b0000000000000000001000: n8470_o = p2;
      22'b0000000000000000000100: n8470_o = p2;
      22'b0000000000000000000010: n8470_o = p2;
      22'b0000000000000000000001: n8470_o = p2;
      default: n8470_o = p2;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8471_o = ie;
      22'b0100000000000000000000: n8471_o = ie;
      22'b0010000000000000000000: n8471_o = ie;
      22'b0001000000000000000000: n8471_o = ie;
      22'b0000100000000000000000: n8471_o = ie;
      22'b0000010000000000000000: n8471_o = s_data;
      22'b0000001000000000000000: n8471_o = ie;
      22'b0000000100000000000000: n8471_o = ie;
      22'b0000000010000000000000: n8471_o = ie;
      22'b0000000001000000000000: n8471_o = ie;
      22'b0000000000100000000000: n8471_o = ie;
      22'b0000000000010000000000: n8471_o = ie;
      22'b0000000000001000000000: n8471_o = ie;
      22'b0000000000000100000000: n8471_o = ie;
      22'b0000000000000010000000: n8471_o = ie;
      22'b0000000000000001000000: n8471_o = ie;
      22'b0000000000000000100000: n8471_o = ie;
      22'b0000000000000000010000: n8471_o = ie;
      22'b0000000000000000001000: n8471_o = ie;
      22'b0000000000000000000100: n8471_o = ie;
      22'b0000000000000000000010: n8471_o = ie;
      22'b0000000000000000000001: n8471_o = ie;
      default: n8471_o = ie;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8472_o = p3;
      22'b0100000000000000000000: n8472_o = p3;
      22'b0010000000000000000000: n8472_o = p3;
      22'b0001000000000000000000: n8472_o = p3;
      22'b0000100000000000000000: n8472_o = s_data;
      22'b0000010000000000000000: n8472_o = p3;
      22'b0000001000000000000000: n8472_o = p3;
      22'b0000000100000000000000: n8472_o = p3;
      22'b0000000010000000000000: n8472_o = p3;
      22'b0000000001000000000000: n8472_o = p3;
      22'b0000000000100000000000: n8472_o = p3;
      22'b0000000000010000000000: n8472_o = p3;
      22'b0000000000001000000000: n8472_o = p3;
      22'b0000000000000100000000: n8472_o = p3;
      22'b0000000000000010000000: n8472_o = p3;
      22'b0000000000000001000000: n8472_o = p3;
      22'b0000000000000000100000: n8472_o = p3;
      22'b0000000000000000010000: n8472_o = p3;
      22'b0000000000000000001000: n8472_o = p3;
      22'b0000000000000000000100: n8472_o = p3;
      22'b0000000000000000000010: n8472_o = p3;
      22'b0000000000000000000001: n8472_o = p3;
      default: n8472_o = p3;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8473_o = ip;
      22'b0100000000000000000000: n8473_o = ip;
      22'b0010000000000000000000: n8473_o = ip;
      22'b0001000000000000000000: n8473_o = s_data;
      22'b0000100000000000000000: n8473_o = ip;
      22'b0000010000000000000000: n8473_o = ip;
      22'b0000001000000000000000: n8473_o = ip;
      22'b0000000100000000000000: n8473_o = ip;
      22'b0000000010000000000000: n8473_o = ip;
      22'b0000000001000000000000: n8473_o = ip;
      22'b0000000000100000000000: n8473_o = ip;
      22'b0000000000010000000000: n8473_o = ip;
      22'b0000000000001000000000: n8473_o = ip;
      22'b0000000000000100000000: n8473_o = ip;
      22'b0000000000000010000000: n8473_o = ip;
      22'b0000000000000001000000: n8473_o = ip;
      22'b0000000000000000100000: n8473_o = ip;
      22'b0000000000000000010000: n8473_o = ip;
      22'b0000000000000000001000: n8473_o = ip;
      22'b0000000000000000000100: n8473_o = ip;
      22'b0000000000000000000010: n8473_o = ip;
      22'b0000000000000000000001: n8473_o = ip;
      default: n8473_o = ip;
    endcase
  assign n8474_o = psw[7:1];
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8475_o = n8474_o;
      22'b0100000000000000000000: n8475_o = n8474_o;
      22'b0010000000000000000000: n8475_o = n8430_o;
      22'b0001000000000000000000: n8475_o = n8474_o;
      22'b0000100000000000000000: n8475_o = n8474_o;
      22'b0000010000000000000000: n8475_o = n8474_o;
      22'b0000001000000000000000: n8475_o = n8474_o;
      22'b0000000100000000000000: n8475_o = n8474_o;
      22'b0000000010000000000000: n8475_o = n8474_o;
      22'b0000000001000000000000: n8475_o = n8474_o;
      22'b0000000000100000000000: n8475_o = n8474_o;
      22'b0000000000010000000000: n8475_o = n8474_o;
      22'b0000000000001000000000: n8475_o = n8474_o;
      22'b0000000000000100000000: n8475_o = n8474_o;
      22'b0000000000000010000000: n8475_o = n8474_o;
      22'b0000000000000001000000: n8475_o = n8474_o;
      22'b0000000000000000100000: n8475_o = n8474_o;
      22'b0000000000000000010000: n8475_o = n8474_o;
      22'b0000000000000000001000: n8475_o = n8474_o;
      22'b0000000000000000000100: n8475_o = n8474_o;
      22'b0000000000000000000010: n8475_o = n8474_o;
      22'b0000000000000000000001: n8475_o = n8474_o;
      default: n8475_o = n8474_o;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8476_o = acc;
      22'b0100000000000000000000: n8476_o = s_data;
      22'b0010000000000000000000: n8476_o = acc;
      22'b0001000000000000000000: n8476_o = acc;
      22'b0000100000000000000000: n8476_o = acc;
      22'b0000010000000000000000: n8476_o = acc;
      22'b0000001000000000000000: n8476_o = acc;
      22'b0000000100000000000000: n8476_o = acc;
      22'b0000000010000000000000: n8476_o = acc;
      22'b0000000001000000000000: n8476_o = acc;
      22'b0000000000100000000000: n8476_o = acc;
      22'b0000000000010000000000: n8476_o = acc;
      22'b0000000000001000000000: n8476_o = acc;
      22'b0000000000000100000000: n8476_o = acc;
      22'b0000000000000010000000: n8476_o = acc;
      22'b0000000000000001000000: n8476_o = acc;
      22'b0000000000000000100000: n8476_o = acc;
      22'b0000000000000000010000: n8476_o = acc;
      22'b0000000000000000001000: n8476_o = acc;
      22'b0000000000000000000100: n8476_o = acc;
      22'b0000000000000000000010: n8476_o = acc;
      22'b0000000000000000000001: n8476_o = acc;
      default: n8476_o = acc;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8477_o = s_data;
      22'b0100000000000000000000: n8477_o = b;
      22'b0010000000000000000000: n8477_o = b;
      22'b0001000000000000000000: n8477_o = b;
      22'b0000100000000000000000: n8477_o = b;
      22'b0000010000000000000000: n8477_o = b;
      22'b0000001000000000000000: n8477_o = b;
      22'b0000000100000000000000: n8477_o = b;
      22'b0000000010000000000000: n8477_o = b;
      22'b0000000001000000000000: n8477_o = b;
      22'b0000000000100000000000: n8477_o = b;
      22'b0000000000010000000000: n8477_o = b;
      22'b0000000000001000000000: n8477_o = b;
      22'b0000000000000100000000: n8477_o = b;
      22'b0000000000000010000000: n8477_o = b;
      22'b0000000000000001000000: n8477_o = b;
      22'b0000000000000000100000: n8477_o = b;
      22'b0000000000000000010000: n8477_o = b;
      22'b0000000000000000001000: n8477_o = b;
      22'b0000000000000000000100: n8477_o = b;
      22'b0000000000000000000010: n8477_o = b;
      22'b0000000000000000000001: n8477_o = b;
      default: n8477_o = b;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8478_o = tsel;
      22'b0100000000000000000000: n8478_o = tsel;
      22'b0010000000000000000000: n8478_o = tsel;
      22'b0001000000000000000000: n8478_o = tsel;
      22'b0000100000000000000000: n8478_o = tsel;
      22'b0000010000000000000000: n8478_o = tsel;
      22'b0000001000000000000000: n8478_o = tsel;
      22'b0000000100000000000000: n8478_o = tsel;
      22'b0000000010000000000000: n8478_o = tsel;
      22'b0000000001000000000000: n8478_o = tsel;
      22'b0000000000100000000000: n8478_o = tsel;
      22'b0000000000010000000000: n8478_o = s_data;
      22'b0000000000001000000000: n8478_o = tsel;
      22'b0000000000000100000000: n8478_o = tsel;
      22'b0000000000000010000000: n8478_o = tsel;
      22'b0000000000000001000000: n8478_o = tsel;
      22'b0000000000000000100000: n8478_o = tsel;
      22'b0000000000000000010000: n8478_o = tsel;
      22'b0000000000000000001000: n8478_o = tsel;
      22'b0000000000000000000100: n8478_o = tsel;
      22'b0000000000000000000010: n8478_o = tsel;
      22'b0000000000000000000001: n8478_o = tsel;
      default: n8478_o = tsel;
    endcase
  /* control_mem_rtl.vhd:1015:15  */
  always @*
    case (n8437_o)
      22'b1000000000000000000000: n8479_o = ssel;
      22'b0100000000000000000000: n8479_o = ssel;
      22'b0010000000000000000000: n8479_o = ssel;
      22'b0001000000000000000000: n8479_o = ssel;
      22'b0000100000000000000000: n8479_o = ssel;
      22'b0000010000000000000000: n8479_o = ssel;
      22'b0000001000000000000000: n8479_o = ssel;
      22'b0000000100000000000000: n8479_o = s_data;
      22'b0000000010000000000000: n8479_o = ssel;
      22'b0000000001000000000000: n8479_o = ssel;
      22'b0000000000100000000000: n8479_o = ssel;
      22'b0000000000010000000000: n8479_o = ssel;
      22'b0000000000001000000000: n8479_o = ssel;
      22'b0000000000000100000000: n8479_o = ssel;
      22'b0000000000000010000000: n8479_o = ssel;
      22'b0000000000000001000000: n8479_o = ssel;
      22'b0000000000000000100000: n8479_o = ssel;
      22'b0000000000000000010000: n8479_o = ssel;
      22'b0000000000000000001000: n8479_o = ssel;
      22'b0000000000000000000100: n8479_o = ssel;
      22'b0000000000000000000010: n8479_o = ssel;
      22'b0000000000000000000001: n8479_o = ssel;
      default: n8479_o = ssel;
    endcase
  /* control_mem_rtl.vhd:1058:46  */
  assign n8480_o = s_adr[7:4];
  /* control_mem_rtl.vhd:1058:61  */
  assign n8482_o = n8480_o == 4'b0010;
  /* control_mem_rtl.vhd:1059:40  */
  assign n8483_o = s_adr[3:0];
  /* control_mem_rtl.vhd:1060:49  */
  assign n8488_o = s_adr == 8'b00000000;
  /* control_mem_rtl.vhd:1062:49  */
  assign n8490_o = s_adr == 8'b00000001;
  /* control_mem_rtl.vhd:1064:49  */
  assign n8492_o = s_adr == 8'b00001000;
  /* control_mem_rtl.vhd:1066:49  */
  assign n8494_o = s_adr == 8'b00001001;
  /* control_mem_rtl.vhd:1068:49  */
  assign n8496_o = s_adr == 8'b00010000;
  /* control_mem_rtl.vhd:1070:49  */
  assign n8498_o = s_adr == 8'b00010001;
  /* control_mem_rtl.vhd:1072:49  */
  assign n8500_o = s_adr == 8'b00011000;
  /* control_mem_rtl.vhd:1074:49  */
  assign n8502_o = s_adr == 8'b00011001;
  /* control_mem_rtl.vhd:1074:13  */
  assign n8503_o = n8502_o ? s_data : s_r1_b3;
  /* control_mem_rtl.vhd:1072:13  */
  assign n8504_o = n8500_o ? s_data : s_r0_b3;
  /* control_mem_rtl.vhd:1072:13  */
  assign n8505_o = n8500_o ? s_r1_b3 : n8503_o;
  /* control_mem_rtl.vhd:1070:13  */
  assign n8506_o = n8498_o ? s_data : s_r1_b2;
  /* control_mem_rtl.vhd:1070:13  */
  assign n8507_o = n8498_o ? s_r0_b3 : n8504_o;
  /* control_mem_rtl.vhd:1070:13  */
  assign n8508_o = n8498_o ? s_r1_b3 : n8505_o;
  /* control_mem_rtl.vhd:1068:13  */
  assign n8509_o = n8496_o ? s_data : s_r0_b2;
  /* control_mem_rtl.vhd:1068:13  */
  assign n8510_o = n8496_o ? s_r1_b2 : n8506_o;
  /* control_mem_rtl.vhd:1068:13  */
  assign n8511_o = n8496_o ? s_r0_b3 : n8507_o;
  /* control_mem_rtl.vhd:1068:13  */
  assign n8512_o = n8496_o ? s_r1_b3 : n8508_o;
  /* control_mem_rtl.vhd:1066:13  */
  assign n8513_o = n8494_o ? s_data : s_r1_b1;
  /* control_mem_rtl.vhd:1066:13  */
  assign n8514_o = n8494_o ? s_r0_b2 : n8509_o;
  /* control_mem_rtl.vhd:1066:13  */
  assign n8515_o = n8494_o ? s_r1_b2 : n8510_o;
  /* control_mem_rtl.vhd:1066:13  */
  assign n8516_o = n8494_o ? s_r0_b3 : n8511_o;
  /* control_mem_rtl.vhd:1066:13  */
  assign n8517_o = n8494_o ? s_r1_b3 : n8512_o;
  /* control_mem_rtl.vhd:1064:13  */
  assign n8518_o = n8492_o ? s_data : s_r0_b1;
  /* control_mem_rtl.vhd:1064:13  */
  assign n8519_o = n8492_o ? s_r1_b1 : n8513_o;
  /* control_mem_rtl.vhd:1064:13  */
  assign n8520_o = n8492_o ? s_r0_b2 : n8514_o;
  /* control_mem_rtl.vhd:1064:13  */
  assign n8521_o = n8492_o ? s_r1_b2 : n8515_o;
  /* control_mem_rtl.vhd:1064:13  */
  assign n8522_o = n8492_o ? s_r0_b3 : n8516_o;
  /* control_mem_rtl.vhd:1064:13  */
  assign n8523_o = n8492_o ? s_r1_b3 : n8517_o;
  /* control_mem_rtl.vhd:1062:13  */
  assign n8524_o = n8490_o ? s_data : s_r1_b0;
  /* control_mem_rtl.vhd:1062:13  */
  assign n8525_o = n8490_o ? s_r0_b1 : n8518_o;
  /* control_mem_rtl.vhd:1062:13  */
  assign n8526_o = n8490_o ? s_r1_b1 : n8519_o;
  /* control_mem_rtl.vhd:1062:13  */
  assign n8527_o = n8490_o ? s_r0_b2 : n8520_o;
  /* control_mem_rtl.vhd:1062:13  */
  assign n8528_o = n8490_o ? s_r1_b2 : n8521_o;
  /* control_mem_rtl.vhd:1062:13  */
  assign n8529_o = n8490_o ? s_r0_b3 : n8522_o;
  /* control_mem_rtl.vhd:1062:13  */
  assign n8530_o = n8490_o ? s_r1_b3 : n8523_o;
  /* control_mem_rtl.vhd:1060:13  */
  assign n8531_o = n8488_o ? s_data : s_r0_b0;
  /* control_mem_rtl.vhd:1060:13  */
  assign n8532_o = n8488_o ? s_r1_b0 : n8524_o;
  /* control_mem_rtl.vhd:1060:13  */
  assign n8533_o = n8488_o ? s_r0_b1 : n8525_o;
  /* control_mem_rtl.vhd:1060:13  */
  assign n8534_o = n8488_o ? s_r1_b1 : n8526_o;
  /* control_mem_rtl.vhd:1060:13  */
  assign n8535_o = n8488_o ? s_r0_b2 : n8527_o;
  /* control_mem_rtl.vhd:1060:13  */
  assign n8536_o = n8488_o ? s_r1_b2 : n8528_o;
  /* control_mem_rtl.vhd:1060:13  */
  assign n8537_o = n8488_o ? s_r0_b3 : n8529_o;
  /* control_mem_rtl.vhd:1060:13  */
  assign n8538_o = n8488_o ? s_r1_b3 : n8530_o;
  /* control_mem_rtl.vhd:1058:13  */
  assign n8539_o = n8482_o ? n9607_o : gprbit;
  /* control_mem_rtl.vhd:1058:13  */
  assign n8540_o = n8482_o ? s_r0_b0 : n8531_o;
  /* control_mem_rtl.vhd:1058:13  */
  assign n8541_o = n8482_o ? s_r1_b0 : n8532_o;
  /* control_mem_rtl.vhd:1058:13  */
  assign n8542_o = n8482_o ? s_r0_b1 : n8533_o;
  /* control_mem_rtl.vhd:1058:13  */
  assign n8543_o = n8482_o ? s_r1_b1 : n8534_o;
  /* control_mem_rtl.vhd:1058:13  */
  assign n8544_o = n8482_o ? s_r0_b2 : n8535_o;
  /* control_mem_rtl.vhd:1058:13  */
  assign n8545_o = n8482_o ? s_r1_b2 : n8536_o;
  /* control_mem_rtl.vhd:1058:13  */
  assign n8546_o = n8482_o ? s_r0_b3 : n8537_o;
  /* control_mem_rtl.vhd:1058:13  */
  assign n8547_o = n8482_o ? s_r1_b3 : n8538_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8549_o = n8388_o ? n8440_o : 1'b0;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8551_o = n8388_o ? n8446_o : 1'b0;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8552_o = n8388_o ? gprbit : n8539_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8553_o = n8388_o ? s_r0_b0 : n8540_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8554_o = n8388_o ? s_r1_b0 : n8541_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8555_o = n8388_o ? s_r0_b1 : n8542_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8556_o = n8388_o ? s_r1_b1 : n8543_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8557_o = n8388_o ? s_r0_b2 : n8544_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8558_o = n8388_o ? s_r1_b2 : n8545_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8559_o = n8388_o ? s_r0_b3 : n8546_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8560_o = n8388_o ? s_r1_b3 : n8547_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8561_o = n8388_o ? n8447_o : s_smodreg;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8562_o = n8388_o ? n8448_o : s_reload;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8563_o = n8388_o ? n8453_o : s_wt;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8564_o = n8388_o ? n8454_o : p0;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8565_o = n8388_o ? n8455_o : dpl;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8566_o = n8388_o ? n8456_o : dph;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8567_o = n8388_o ? n8457_o : pcon;
  assign n8568_o = tcon[0];
  assign n8569_o = tcon[2];
  assign n8570_o = tcon[4];
  assign n8571_o = tcon[6];
  assign n8572_o = {n8320_o, n8571_o, n8318_o, n8570_o, n8304_o, n8569_o, n8316_o, n8568_o};
  /* control_mem_rtl.vhd:1014:13  */
  assign n8573_o = n8388_o ? n8463_o : n8572_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8574_o = n8388_o ? n8464_o : tmod;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8575_o = n8388_o ? n8465_o : p1;
  assign n8576_o = scon[7:2];
  assign n8577_o = {n8576_o, n8324_o, n8322_o};
  /* control_mem_rtl.vhd:1014:13  */
  assign n8578_o = n8388_o ? n8468_o : n8577_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8579_o = n8388_o ? n8469_o : sbuf;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8580_o = n8388_o ? n8470_o : p2;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8581_o = n8388_o ? n8471_o : ie;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8582_o = n8388_o ? n8472_o : p3;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8583_o = n8388_o ? n8473_o : ip;
  assign n8584_o = psw[7:1];
  /* control_mem_rtl.vhd:1014:13  */
  assign n8585_o = n8388_o ? n8475_o : n8584_o;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8586_o = n8388_o ? n8476_o : acc;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8587_o = n8388_o ? n8477_o : b;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8588_o = n8388_o ? n8478_o : tsel;
  /* control_mem_rtl.vhd:1014:13  */
  assign n8589_o = n8388_o ? n8479_o : ssel;
  /* control_mem_rtl.vhd:991:11  */
  assign n8591_o = s_regs_wr_en == 3'b100;
  /* control_mem_rtl.vhd:991:22  */
  assign n8593_o = s_regs_wr_en == 3'b101;
  /* control_mem_rtl.vhd:991:22  */
  assign n8594_o = n8591_o | n8593_o;
  /* control_mem_rtl.vhd:1080:27  */
  assign n8595_o = ~s_intblock;
  /* control_mem_rtl.vhd:1080:32  */
  assign n8596_o = n8595_o & s_intpre;
  /* control_mem_rtl.vhd:1080:58  */
  assign n8598_o = state == 3'b001;
  /* control_mem_rtl.vhd:1080:49  */
  assign n8599_o = n8596_o & n8598_o;
  /* control_mem_rtl.vhd:1080:66  */
  assign n8600_o = n8599_o | s_intpre2;
  /* control_mem_rtl.vhd:1081:27  */
  assign n8602_o = s_command != 8'b10000010;
  /* control_mem_rtl.vhd:1082:27  */
  assign n8604_o = s_command != 8'b10110000;
  /* control_mem_rtl.vhd:1081:40  */
  assign n8605_o = n8602_o & n8604_o;
  /* control_mem_rtl.vhd:1083:27  */
  assign n8607_o = s_command != 8'b10100010;
  /* control_mem_rtl.vhd:1082:41  */
  assign n8608_o = n8605_o & n8607_o;
  /* control_mem_rtl.vhd:1084:27  */
  assign n8610_o = s_command != 8'b01110010;
  /* control_mem_rtl.vhd:1083:40  */
  assign n8611_o = n8608_o & n8610_o;
  /* control_mem_rtl.vhd:1085:27  */
  assign n8613_o = s_command != 8'b10100000;
  /* control_mem_rtl.vhd:1084:40  */
  assign n8614_o = n8611_o & n8613_o;
  /* control_mem_rtl.vhd:1080:83  */
  assign n8615_o = n8600_o | n8614_o;
  /* control_mem_rtl.vhd:1086:23  */
  assign n8616_o = s_adr[7];
  /* control_mem_rtl.vhd:1087:27  */
  assign n8617_o = s_adr[6:3];
  /* control_mem_rtl.vhd:1089:42  */
  assign n8618_o = s_adr[2:0];
  /* control_mem_rtl.vhd:1088:19  */
  assign n8623_o = n8617_o == 4'b0000;
  /* control_mem_rtl.vhd:1091:52  */
  assign n8624_o = s_adr[2:0];
  assign n8627_o = tcon[0];
  assign n8628_o = tcon[2];
  assign n8629_o = tcon[4];
  assign n8630_o = tcon[6];
  assign n8631_o = {n8320_o, n8630_o, n8318_o, n8629_o, n8304_o, n8628_o, n8316_o, n8627_o};
  /* control_mem_rtl.vhd:1090:19  */
  assign n8634_o = n8617_o == 4'b0001;
  /* control_mem_rtl.vhd:1093:42  */
  assign n8635_o = s_adr[2:0];
  /* control_mem_rtl.vhd:1092:19  */
  assign n8640_o = n8617_o == 4'b0010;
  /* control_mem_rtl.vhd:1095:52  */
  assign n8641_o = s_adr[2:0];
  assign n8644_o = scon[7:2];
  assign n8645_o = {n8644_o, n8324_o, n8322_o};
  /* control_mem_rtl.vhd:1094:19  */
  assign n8648_o = n8617_o == 4'b0011;
  /* control_mem_rtl.vhd:1097:42  */
  assign n8649_o = s_adr[2:0];
  /* control_mem_rtl.vhd:1096:19  */
  assign n8654_o = n8617_o == 4'b0100;
  /* control_mem_rtl.vhd:1099:42  */
  assign n8655_o = s_adr[2:0];
  /* control_mem_rtl.vhd:1098:19  */
  assign n8660_o = n8617_o == 4'b0101;
  /* control_mem_rtl.vhd:1101:42  */
  assign n8661_o = s_adr[2:0];
  /* control_mem_rtl.vhd:1100:19  */
  assign n8666_o = n8617_o == 4'b0110;
  /* control_mem_rtl.vhd:1103:42  */
  assign n8667_o = s_adr[2:0];
  /* control_mem_rtl.vhd:1102:19  */
  assign n8672_o = n8617_o == 4'b0111;
  /* control_mem_rtl.vhd:1105:31  */
  assign n8673_o = s_adr[2:0];
  /* control_mem_rtl.vhd:1106:23  */
  assign n8675_o = n8673_o == 3'b000;
  /* control_mem_rtl.vhd:1107:23  */
  assign n8677_o = n8673_o == 3'b001;
  /* control_mem_rtl.vhd:1108:23  */
  assign n8679_o = n8673_o == 3'b010;
  /* control_mem_rtl.vhd:1109:23  */
  assign n8681_o = n8673_o == 3'b011;
  /* control_mem_rtl.vhd:1110:23  */
  assign n8683_o = n8673_o == 3'b100;
  /* control_mem_rtl.vhd:1111:23  */
  assign n8685_o = n8673_o == 3'b101;
  /* control_mem_rtl.vhd:1112:23  */
  assign n8687_o = n8673_o == 3'b110;
  /* control_mem_rtl.vhd:1113:23  */
  assign n8689_o = n8673_o == 3'b111;
  assign n8690_o = {n8689_o, n8687_o, n8685_o, n8683_o, n8681_o, n8679_o, n8677_o, n8675_o};
  assign n8691_o = psw[1];
  /* control_mem_rtl.vhd:1105:21  */
  always @*
    case (n8690_o)
      8'b10000000: n8692_o = n8691_o;
      8'b01000000: n8692_o = n8691_o;
      8'b00100000: n8692_o = n8691_o;
      8'b00010000: n8692_o = n8691_o;
      8'b00001000: n8692_o = n8691_o;
      8'b00000100: n8692_o = n8691_o;
      8'b00000010: n8692_o = s_bdata;
      8'b00000001: n8692_o = n8691_o;
      default: n8692_o = n8691_o;
    endcase
  assign n8693_o = psw[2];
  /* control_mem_rtl.vhd:1105:21  */
  always @*
    case (n8690_o)
      8'b10000000: n8694_o = n8693_o;
      8'b01000000: n8694_o = n8693_o;
      8'b00100000: n8694_o = n8693_o;
      8'b00010000: n8694_o = n8693_o;
      8'b00001000: n8694_o = n8693_o;
      8'b00000100: n8694_o = s_bdata;
      8'b00000010: n8694_o = n8693_o;
      8'b00000001: n8694_o = n8693_o;
      default: n8694_o = n8693_o;
    endcase
  assign n8695_o = psw[3];
  /* control_mem_rtl.vhd:1105:21  */
  always @*
    case (n8690_o)
      8'b10000000: n8696_o = n8695_o;
      8'b01000000: n8696_o = n8695_o;
      8'b00100000: n8696_o = n8695_o;
      8'b00010000: n8696_o = n8695_o;
      8'b00001000: n8696_o = s_bdata;
      8'b00000100: n8696_o = n8695_o;
      8'b00000010: n8696_o = n8695_o;
      8'b00000001: n8696_o = n8695_o;
      default: n8696_o = n8695_o;
    endcase
  assign n8697_o = psw[4];
  /* control_mem_rtl.vhd:1105:21  */
  always @*
    case (n8690_o)
      8'b10000000: n8698_o = n8697_o;
      8'b01000000: n8698_o = n8697_o;
      8'b00100000: n8698_o = n8697_o;
      8'b00010000: n8698_o = s_bdata;
      8'b00001000: n8698_o = n8697_o;
      8'b00000100: n8698_o = n8697_o;
      8'b00000010: n8698_o = n8697_o;
      8'b00000001: n8698_o = n8697_o;
      default: n8698_o = n8697_o;
    endcase
  assign n8699_o = psw[5];
  /* control_mem_rtl.vhd:1105:21  */
  always @*
    case (n8690_o)
      8'b10000000: n8700_o = n8699_o;
      8'b01000000: n8700_o = n8699_o;
      8'b00100000: n8700_o = s_bdata;
      8'b00010000: n8700_o = n8699_o;
      8'b00001000: n8700_o = n8699_o;
      8'b00000100: n8700_o = n8699_o;
      8'b00000010: n8700_o = n8699_o;
      8'b00000001: n8700_o = n8699_o;
      default: n8700_o = n8699_o;
    endcase
  assign n8701_o = psw[6];
  /* control_mem_rtl.vhd:1105:21  */
  always @*
    case (n8690_o)
      8'b10000000: n8702_o = n8701_o;
      8'b01000000: n8702_o = s_bdata;
      8'b00100000: n8702_o = n8701_o;
      8'b00010000: n8702_o = n8701_o;
      8'b00001000: n8702_o = n8701_o;
      8'b00000100: n8702_o = n8701_o;
      8'b00000010: n8702_o = n8701_o;
      8'b00000001: n8702_o = n8701_o;
      default: n8702_o = n8701_o;
    endcase
  assign n8703_o = psw[7];
  /* control_mem_rtl.vhd:1105:21  */
  always @*
    case (n8690_o)
      8'b10000000: n8704_o = s_bdata;
      8'b01000000: n8704_o = n8703_o;
      8'b00100000: n8704_o = n8703_o;
      8'b00010000: n8704_o = n8703_o;
      8'b00001000: n8704_o = n8703_o;
      8'b00000100: n8704_o = n8703_o;
      8'b00000010: n8704_o = n8703_o;
      8'b00000001: n8704_o = n8703_o;
      default: n8704_o = n8703_o;
    endcase
  /* control_mem_rtl.vhd:1104:19  */
  assign n8706_o = n8617_o == 4'b1010;
  /* control_mem_rtl.vhd:1117:43  */
  assign n8707_o = s_adr[2:0];
  /* control_mem_rtl.vhd:1116:19  */
  assign n8712_o = n8617_o == 4'b1100;
  /* control_mem_rtl.vhd:1119:41  */
  assign n8713_o = s_adr[2:0];
  /* control_mem_rtl.vhd:1118:19  */
  assign n8718_o = n8617_o == 4'b1110;
  assign n8719_o = {n8718_o, n8712_o, n8706_o, n8672_o, n8666_o, n8660_o, n8654_o, n8648_o, n8640_o, n8634_o, n8623_o};
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8720_o = p0;
      11'b01000000000: n8720_o = p0;
      11'b00100000000: n8720_o = p0;
      11'b00010000000: n8720_o = p0;
      11'b00001000000: n8720_o = p0;
      11'b00000100000: n8720_o = p0;
      11'b00000010000: n8720_o = p0;
      11'b00000001000: n8720_o = p0;
      11'b00000000100: n8720_o = p0;
      11'b00000000010: n8720_o = p0;
      11'b00000000001: n8720_o = n9642_o;
      default: n8720_o = p0;
    endcase
  assign n8721_o = tcon[0];
  assign n8722_o = tcon[2];
  assign n8723_o = tcon[4];
  assign n8724_o = tcon[6];
  assign n8725_o = {n8320_o, n8724_o, n8318_o, n8723_o, n8304_o, n8722_o, n8316_o, n8721_o};
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8726_o = n8725_o;
      11'b01000000000: n8726_o = n8725_o;
      11'b00100000000: n8726_o = n8725_o;
      11'b00010000000: n8726_o = n8725_o;
      11'b00001000000: n8726_o = n8725_o;
      11'b00000100000: n8726_o = n8725_o;
      11'b00000010000: n8726_o = n8725_o;
      11'b00000001000: n8726_o = n8725_o;
      11'b00000000100: n8726_o = n8725_o;
      11'b00000000010: n8726_o = n9677_o;
      11'b00000000001: n8726_o = n8725_o;
      default: n8726_o = n8725_o;
    endcase
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8727_o = p1;
      11'b01000000000: n8727_o = p1;
      11'b00100000000: n8727_o = p1;
      11'b00010000000: n8727_o = p1;
      11'b00001000000: n8727_o = p1;
      11'b00000100000: n8727_o = p1;
      11'b00000010000: n8727_o = p1;
      11'b00000001000: n8727_o = p1;
      11'b00000000100: n8727_o = n9712_o;
      11'b00000000010: n8727_o = p1;
      11'b00000000001: n8727_o = p1;
      default: n8727_o = p1;
    endcase
  assign n8728_o = scon[7:2];
  assign n8729_o = {n8728_o, n8324_o, n8322_o};
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8730_o = n8729_o;
      11'b01000000000: n8730_o = n8729_o;
      11'b00100000000: n8730_o = n8729_o;
      11'b00010000000: n8730_o = n8729_o;
      11'b00001000000: n8730_o = n8729_o;
      11'b00000100000: n8730_o = n8729_o;
      11'b00000010000: n8730_o = n8729_o;
      11'b00000001000: n8730_o = n9747_o;
      11'b00000000100: n8730_o = n8729_o;
      11'b00000000010: n8730_o = n8729_o;
      11'b00000000001: n8730_o = n8729_o;
      default: n8730_o = n8729_o;
    endcase
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8731_o = p2;
      11'b01000000000: n8731_o = p2;
      11'b00100000000: n8731_o = p2;
      11'b00010000000: n8731_o = p2;
      11'b00001000000: n8731_o = p2;
      11'b00000100000: n8731_o = p2;
      11'b00000010000: n8731_o = n9782_o;
      11'b00000001000: n8731_o = p2;
      11'b00000000100: n8731_o = p2;
      11'b00000000010: n8731_o = p2;
      11'b00000000001: n8731_o = p2;
      default: n8731_o = p2;
    endcase
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8732_o = ie;
      11'b01000000000: n8732_o = ie;
      11'b00100000000: n8732_o = ie;
      11'b00010000000: n8732_o = ie;
      11'b00001000000: n8732_o = ie;
      11'b00000100000: n8732_o = n9817_o;
      11'b00000010000: n8732_o = ie;
      11'b00000001000: n8732_o = ie;
      11'b00000000100: n8732_o = ie;
      11'b00000000010: n8732_o = ie;
      11'b00000000001: n8732_o = ie;
      default: n8732_o = ie;
    endcase
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8733_o = p3;
      11'b01000000000: n8733_o = p3;
      11'b00100000000: n8733_o = p3;
      11'b00010000000: n8733_o = p3;
      11'b00001000000: n8733_o = n9852_o;
      11'b00000100000: n8733_o = p3;
      11'b00000010000: n8733_o = p3;
      11'b00000001000: n8733_o = p3;
      11'b00000000100: n8733_o = p3;
      11'b00000000010: n8733_o = p3;
      11'b00000000001: n8733_o = p3;
      default: n8733_o = p3;
    endcase
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8734_o = ip;
      11'b01000000000: n8734_o = ip;
      11'b00100000000: n8734_o = ip;
      11'b00010000000: n8734_o = n9887_o;
      11'b00001000000: n8734_o = ip;
      11'b00000100000: n8734_o = ip;
      11'b00000010000: n8734_o = ip;
      11'b00000001000: n8734_o = ip;
      11'b00000000100: n8734_o = ip;
      11'b00000000010: n8734_o = ip;
      11'b00000000001: n8734_o = ip;
      default: n8734_o = ip;
    endcase
  assign n8735_o = psw[1];
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8736_o = n8735_o;
      11'b01000000000: n8736_o = n8735_o;
      11'b00100000000: n8736_o = n8692_o;
      11'b00010000000: n8736_o = n8735_o;
      11'b00001000000: n8736_o = n8735_o;
      11'b00000100000: n8736_o = n8735_o;
      11'b00000010000: n8736_o = n8735_o;
      11'b00000001000: n8736_o = n8735_o;
      11'b00000000100: n8736_o = n8735_o;
      11'b00000000010: n8736_o = n8735_o;
      11'b00000000001: n8736_o = n8735_o;
      default: n8736_o = n8735_o;
    endcase
  assign n8737_o = psw[2];
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8738_o = n8737_o;
      11'b01000000000: n8738_o = n8737_o;
      11'b00100000000: n8738_o = n8694_o;
      11'b00010000000: n8738_o = n8737_o;
      11'b00001000000: n8738_o = n8737_o;
      11'b00000100000: n8738_o = n8737_o;
      11'b00000010000: n8738_o = n8737_o;
      11'b00000001000: n8738_o = n8737_o;
      11'b00000000100: n8738_o = n8737_o;
      11'b00000000010: n8738_o = n8737_o;
      11'b00000000001: n8738_o = n8737_o;
      default: n8738_o = n8737_o;
    endcase
  assign n8739_o = psw[3];
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8740_o = n8739_o;
      11'b01000000000: n8740_o = n8739_o;
      11'b00100000000: n8740_o = n8696_o;
      11'b00010000000: n8740_o = n8739_o;
      11'b00001000000: n8740_o = n8739_o;
      11'b00000100000: n8740_o = n8739_o;
      11'b00000010000: n8740_o = n8739_o;
      11'b00000001000: n8740_o = n8739_o;
      11'b00000000100: n8740_o = n8739_o;
      11'b00000000010: n8740_o = n8739_o;
      11'b00000000001: n8740_o = n8739_o;
      default: n8740_o = n8739_o;
    endcase
  assign n8741_o = psw[4];
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8742_o = n8741_o;
      11'b01000000000: n8742_o = n8741_o;
      11'b00100000000: n8742_o = n8698_o;
      11'b00010000000: n8742_o = n8741_o;
      11'b00001000000: n8742_o = n8741_o;
      11'b00000100000: n8742_o = n8741_o;
      11'b00000010000: n8742_o = n8741_o;
      11'b00000001000: n8742_o = n8741_o;
      11'b00000000100: n8742_o = n8741_o;
      11'b00000000010: n8742_o = n8741_o;
      11'b00000000001: n8742_o = n8741_o;
      default: n8742_o = n8741_o;
    endcase
  assign n8743_o = psw[5];
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8744_o = n8743_o;
      11'b01000000000: n8744_o = n8743_o;
      11'b00100000000: n8744_o = n8700_o;
      11'b00010000000: n8744_o = n8743_o;
      11'b00001000000: n8744_o = n8743_o;
      11'b00000100000: n8744_o = n8743_o;
      11'b00000010000: n8744_o = n8743_o;
      11'b00000001000: n8744_o = n8743_o;
      11'b00000000100: n8744_o = n8743_o;
      11'b00000000010: n8744_o = n8743_o;
      11'b00000000001: n8744_o = n8743_o;
      default: n8744_o = n8743_o;
    endcase
  assign n8745_o = psw[6];
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8746_o = n8745_o;
      11'b01000000000: n8746_o = n8745_o;
      11'b00100000000: n8746_o = n8702_o;
      11'b00010000000: n8746_o = n8745_o;
      11'b00001000000: n8746_o = n8745_o;
      11'b00000100000: n8746_o = n8745_o;
      11'b00000010000: n8746_o = n8745_o;
      11'b00000001000: n8746_o = n8745_o;
      11'b00000000100: n8746_o = n8745_o;
      11'b00000000010: n8746_o = n8745_o;
      11'b00000000001: n8746_o = n8745_o;
      default: n8746_o = n8745_o;
    endcase
  assign n8747_o = psw[7];
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8748_o = n8747_o;
      11'b01000000000: n8748_o = n8747_o;
      11'b00100000000: n8748_o = n8704_o;
      11'b00010000000: n8748_o = n8747_o;
      11'b00001000000: n8748_o = n8747_o;
      11'b00000100000: n8748_o = n8747_o;
      11'b00000010000: n8748_o = n8747_o;
      11'b00000001000: n8748_o = n8747_o;
      11'b00000000100: n8748_o = n8747_o;
      11'b00000000010: n8748_o = n8747_o;
      11'b00000000001: n8748_o = n8747_o;
      default: n8748_o = n8747_o;
    endcase
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8749_o = acc;
      11'b01000000000: n8749_o = n9922_o;
      11'b00100000000: n8749_o = acc;
      11'b00010000000: n8749_o = acc;
      11'b00001000000: n8749_o = acc;
      11'b00000100000: n8749_o = acc;
      11'b00000010000: n8749_o = acc;
      11'b00000001000: n8749_o = acc;
      11'b00000000100: n8749_o = acc;
      11'b00000000010: n8749_o = acc;
      11'b00000000001: n8749_o = acc;
      default: n8749_o = acc;
    endcase
  /* control_mem_rtl.vhd:1087:17  */
  always @*
    case (n8719_o)
      11'b10000000000: n8750_o = n9957_o;
      11'b01000000000: n8750_o = b;
      11'b00100000000: n8750_o = b;
      11'b00010000000: n8750_o = b;
      11'b00001000000: n8750_o = b;
      11'b00000100000: n8750_o = b;
      11'b00000010000: n8750_o = b;
      11'b00000001000: n8750_o = b;
      11'b00000000100: n8750_o = b;
      11'b00000000010: n8750_o = b;
      11'b00000000001: n8750_o = b;
      default: n8750_o = b;
    endcase
  /* control_mem_rtl.vhd:1123:42  */
  assign n8751_o = s_adr[6:3];
  /* control_mem_rtl.vhd:1124:42  */
  assign n8754_o = s_adr[2:0];
  /* control_mem_rtl.vhd:1086:15  */
  assign n8759_o = n8616_o ? gprbit : n10481_o;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8760_o = n8781_o ? n8720_o : p0;
  assign n8761_o = tcon[0];
  assign n8762_o = tcon[2];
  assign n8763_o = tcon[4];
  assign n8764_o = tcon[6];
  assign n8765_o = {n8320_o, n8764_o, n8318_o, n8763_o, n8304_o, n8762_o, n8316_o, n8761_o};
  /* control_mem_rtl.vhd:1086:15  */
  assign n8766_o = n8616_o ? n8726_o : n8765_o;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8767_o = n8788_o ? n8727_o : p1;
  assign n8768_o = scon[7:2];
  assign n8769_o = {n8768_o, n8324_o, n8322_o};
  /* control_mem_rtl.vhd:1086:15  */
  assign n8770_o = n8616_o ? n8730_o : n8769_o;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8771_o = n8792_o ? n8731_o : p2;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8772_o = n8793_o ? n8732_o : ie;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8773_o = n8794_o ? n8733_o : p3;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8774_o = n8795_o ? n8734_o : ip;
  assign n8775_o = {n8748_o, n8746_o, n8744_o, n8742_o, n8740_o, n8738_o, n8736_o};
  assign n8776_o = psw[7:1];
  /* control_mem_rtl.vhd:1086:15  */
  assign n8777_o = n8616_o ? n8775_o : n8776_o;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8778_o = n8801_o ? n8749_o : acc;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8779_o = n8802_o ? n8750_o : b;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8780_o = n8615_o ? n8759_o : gprbit;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8781_o = n8615_o & n8616_o;
  assign n8782_o = tcon[0];
  assign n8783_o = tcon[2];
  assign n8784_o = tcon[4];
  assign n8785_o = tcon[6];
  assign n8786_o = {n8320_o, n8785_o, n8318_o, n8784_o, n8304_o, n8783_o, n8316_o, n8782_o};
  /* control_mem_rtl.vhd:1080:13  */
  assign n8787_o = n8615_o ? n8766_o : n8786_o;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8788_o = n8615_o & n8616_o;
  assign n8789_o = scon[7:2];
  assign n8790_o = {n8789_o, n8324_o, n8322_o};
  /* control_mem_rtl.vhd:1080:13  */
  assign n8791_o = n8615_o ? n8770_o : n8790_o;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8792_o = n8615_o & n8616_o;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8793_o = n8615_o & n8616_o;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8794_o = n8615_o & n8616_o;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8795_o = n8615_o & n8616_o;
  assign n8796_o = n8777_o[5:0];
  assign n8797_o = psw[6:1];
  /* control_mem_rtl.vhd:1080:13  */
  assign n8798_o = n8615_o ? n8796_o : n8797_o;
  assign n8799_o = n8777_o[6];
  /* control_mem_rtl.vhd:1080:13  */
  assign n8800_o = n8615_o ? n8799_o : s_bdata;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8801_o = n8615_o & n8616_o;
  /* control_mem_rtl.vhd:1080:13  */
  assign n8802_o = n8615_o & n8616_o;
  /* control_mem_rtl.vhd:1079:11  */
  assign n8804_o = s_regs_wr_en == 3'b110;
  /* control_mem_rtl.vhd:1133:35  */
  assign n8805_o = new_cy_i[1];
  /* control_mem_rtl.vhd:1131:15  */
  assign n8807_o = s_command == 8'b11010100;
  /* control_mem_rtl.vhd:1131:25  */
  assign n8809_o = s_command == 8'b00110011;
  /* control_mem_rtl.vhd:1131:25  */
  assign n8810_o = n8807_o | n8809_o;
  /* control_mem_rtl.vhd:1131:33  */
  assign n8812_o = s_command == 8'b00010011;
  /* control_mem_rtl.vhd:1131:33  */
  assign n8813_o = n8810_o | n8812_o;
  /* control_mem_rtl.vhd:1134:15  */
  assign n8816_o = s_command == 8'b10000100;
  /* control_mem_rtl.vhd:1134:27  */
  assign n8818_o = s_command == 8'b10100100;
  /* control_mem_rtl.vhd:1134:27  */
  assign n8819_o = n8816_o | n8818_o;
  assign n8820_o = {n8819_o, n8813_o};
  assign n8821_o = psw[2];
  /* control_mem_rtl.vhd:1130:13  */
  always @*
    case (n8820_o)
      2'b10: n8822_o = new_ov_i;
      2'b01: n8822_o = n8821_o;
      default: n8822_o = n8821_o;
    endcase
  assign n8823_o = psw[7];
  /* control_mem_rtl.vhd:1130:13  */
  always @*
    case (n8820_o)
      2'b10: n8824_o = 1'b0;
      2'b01: n8824_o = n8805_o;
      default: n8824_o = n8823_o;
    endcase
  /* control_mem_rtl.vhd:1130:13  */
  always @*
    case (n8820_o)
      2'b10: n8825_o = s_data;
      2'b01: n8825_o = s_data;
      default: n8825_o = acc;
    endcase
  /* control_mem_rtl.vhd:1130:13  */
  always @*
    case (n8820_o)
      2'b10: n8826_o = aludatb_i;
      2'b01: n8826_o = b;
      default: n8826_o = b;
    endcase
  /* control_mem_rtl.vhd:1129:11  */
  assign n8828_o = s_regs_wr_en == 3'b111;
  assign n8829_o = {n8828_o, n8804_o, n8594_o, n8354_o, n8350_o, n8348_o};
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8831_o = 1'b0;
      6'b010000: n8831_o = 1'b0;
      6'b001000: n8831_o = n8549_o;
      6'b000100: n8831_o = 1'b0;
      6'b000010: n8831_o = 1'b0;
      6'b000001: n8831_o = 1'b0;
      default: n8831_o = 1'b0;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8834_o = 1'b0;
      6'b010000: n8834_o = 1'b0;
      6'b001000: n8834_o = n8551_o;
      6'b000100: n8834_o = 1'b0;
      6'b000010: n8834_o = 1'b0;
      6'b000001: n8834_o = 1'b0;
      default: n8834_o = 1'b0;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8836_o = gprbit;
      6'b010000: n8836_o = n8780_o;
      6'b001000: n8836_o = n8552_o;
      6'b000100: n8836_o = gprbit;
      6'b000010: n8836_o = gprbit;
      6'b000001: n8836_o = gprbit;
      default: n8836_o = gprbit;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8837_o = s_r0_b0;
      6'b010000: n8837_o = s_r0_b0;
      6'b001000: n8837_o = n8553_o;
      6'b000100: n8837_o = s_r0_b0;
      6'b000010: n8837_o = s_r0_b0;
      6'b000001: n8837_o = s_r0_b0;
      default: n8837_o = s_r0_b0;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8838_o = s_r1_b0;
      6'b010000: n8838_o = s_r1_b0;
      6'b001000: n8838_o = n8554_o;
      6'b000100: n8838_o = s_r1_b0;
      6'b000010: n8838_o = s_r1_b0;
      6'b000001: n8838_o = s_r1_b0;
      default: n8838_o = s_r1_b0;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8839_o = s_r0_b1;
      6'b010000: n8839_o = s_r0_b1;
      6'b001000: n8839_o = n8555_o;
      6'b000100: n8839_o = s_r0_b1;
      6'b000010: n8839_o = s_r0_b1;
      6'b000001: n8839_o = s_r0_b1;
      default: n8839_o = s_r0_b1;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8840_o = s_r1_b1;
      6'b010000: n8840_o = s_r1_b1;
      6'b001000: n8840_o = n8556_o;
      6'b000100: n8840_o = s_r1_b1;
      6'b000010: n8840_o = s_r1_b1;
      6'b000001: n8840_o = s_r1_b1;
      default: n8840_o = s_r1_b1;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8841_o = s_r0_b2;
      6'b010000: n8841_o = s_r0_b2;
      6'b001000: n8841_o = n8557_o;
      6'b000100: n8841_o = s_r0_b2;
      6'b000010: n8841_o = s_r0_b2;
      6'b000001: n8841_o = s_r0_b2;
      default: n8841_o = s_r0_b2;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8842_o = s_r1_b2;
      6'b010000: n8842_o = s_r1_b2;
      6'b001000: n8842_o = n8558_o;
      6'b000100: n8842_o = s_r1_b2;
      6'b000010: n8842_o = s_r1_b2;
      6'b000001: n8842_o = s_r1_b2;
      default: n8842_o = s_r1_b2;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8843_o = s_r0_b3;
      6'b010000: n8843_o = s_r0_b3;
      6'b001000: n8843_o = n8559_o;
      6'b000100: n8843_o = s_r0_b3;
      6'b000010: n8843_o = s_r0_b3;
      6'b000001: n8843_o = s_r0_b3;
      default: n8843_o = s_r0_b3;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8844_o = s_r1_b3;
      6'b010000: n8844_o = s_r1_b3;
      6'b001000: n8844_o = n8560_o;
      6'b000100: n8844_o = s_r1_b3;
      6'b000010: n8844_o = s_r1_b3;
      6'b000001: n8844_o = s_r1_b3;
      default: n8844_o = s_r1_b3;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8845_o = s_smodreg;
      6'b010000: n8845_o = s_smodreg;
      6'b001000: n8845_o = n8561_o;
      6'b000100: n8845_o = s_smodreg;
      6'b000010: n8845_o = s_smodreg;
      6'b000001: n8845_o = s_smodreg;
      default: n8845_o = s_smodreg;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8846_o = s_reload;
      6'b010000: n8846_o = s_reload;
      6'b001000: n8846_o = n8562_o;
      6'b000100: n8846_o = s_reload;
      6'b000010: n8846_o = s_reload;
      6'b000001: n8846_o = s_reload;
      default: n8846_o = s_reload;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8847_o = s_wt;
      6'b010000: n8847_o = s_wt;
      6'b001000: n8847_o = n8563_o;
      6'b000100: n8847_o = s_wt;
      6'b000010: n8847_o = s_wt;
      6'b000001: n8847_o = s_wt;
      default: n8847_o = s_wt;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8848_o = p0;
      6'b010000: n8848_o = n8760_o;
      6'b001000: n8848_o = n8564_o;
      6'b000100: n8848_o = p0;
      6'b000010: n8848_o = p0;
      6'b000001: n8848_o = p0;
      default: n8848_o = p0;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8849_o = sp;
      6'b010000: n8849_o = sp;
      6'b001000: n8849_o = n8387_o;
      6'b000100: n8849_o = sp;
      6'b000010: n8849_o = sp;
      6'b000001: n8849_o = n8346_o;
      default: n8849_o = sp;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8850_o = dpl;
      6'b010000: n8850_o = dpl;
      6'b001000: n8850_o = n8565_o;
      6'b000100: n8850_o = dpl;
      6'b000010: n8850_o = dpl;
      6'b000001: n8850_o = dpl;
      default: n8850_o = dpl;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8851_o = dph;
      6'b010000: n8851_o = dph;
      6'b001000: n8851_o = n8566_o;
      6'b000100: n8851_o = dph;
      6'b000010: n8851_o = dph;
      6'b000001: n8851_o = dph;
      default: n8851_o = dph;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8852_o = pcon;
      6'b010000: n8852_o = pcon;
      6'b001000: n8852_o = n8567_o;
      6'b000100: n8852_o = pcon;
      6'b000010: n8852_o = pcon;
      6'b000001: n8852_o = pcon;
      default: n8852_o = pcon;
    endcase
  assign n8853_o = tcon[0];
  assign n8854_o = tcon[2];
  assign n8855_o = tcon[4];
  assign n8856_o = tcon[6];
  assign n8857_o = {n8320_o, n8856_o, n8318_o, n8855_o, n8304_o, n8854_o, n8316_o, n8853_o};
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8858_o = n8857_o;
      6'b010000: n8858_o = n8787_o;
      6'b001000: n8858_o = n8573_o;
      6'b000100: n8858_o = n8857_o;
      6'b000010: n8858_o = n8857_o;
      6'b000001: n8858_o = n8857_o;
      default: n8858_o = n8857_o;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8859_o = tmod;
      6'b010000: n8859_o = tmod;
      6'b001000: n8859_o = n8574_o;
      6'b000100: n8859_o = tmod;
      6'b000010: n8859_o = tmod;
      6'b000001: n8859_o = tmod;
      default: n8859_o = tmod;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8860_o = p1;
      6'b010000: n8860_o = n8767_o;
      6'b001000: n8860_o = n8575_o;
      6'b000100: n8860_o = p1;
      6'b000010: n8860_o = p1;
      6'b000001: n8860_o = p1;
      default: n8860_o = p1;
    endcase
  assign n8861_o = scon[7:2];
  assign n8862_o = {n8861_o, n8324_o, n8322_o};
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8863_o = n8862_o;
      6'b010000: n8863_o = n8791_o;
      6'b001000: n8863_o = n8578_o;
      6'b000100: n8863_o = n8862_o;
      6'b000010: n8863_o = n8862_o;
      6'b000001: n8863_o = n8862_o;
      default: n8863_o = n8862_o;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8864_o = sbuf;
      6'b010000: n8864_o = sbuf;
      6'b001000: n8864_o = n8579_o;
      6'b000100: n8864_o = sbuf;
      6'b000010: n8864_o = sbuf;
      6'b000001: n8864_o = sbuf;
      default: n8864_o = sbuf;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8865_o = p2;
      6'b010000: n8865_o = n8771_o;
      6'b001000: n8865_o = n8580_o;
      6'b000100: n8865_o = p2;
      6'b000010: n8865_o = p2;
      6'b000001: n8865_o = p2;
      default: n8865_o = p2;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8866_o = ie;
      6'b010000: n8866_o = n8772_o;
      6'b001000: n8866_o = n8581_o;
      6'b000100: n8866_o = ie;
      6'b000010: n8866_o = ie;
      6'b000001: n8866_o = ie;
      default: n8866_o = ie;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8867_o = p3;
      6'b010000: n8867_o = n8773_o;
      6'b001000: n8867_o = n8582_o;
      6'b000100: n8867_o = p3;
      6'b000010: n8867_o = p3;
      6'b000001: n8867_o = p3;
      default: n8867_o = p3;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8868_o = ip;
      6'b010000: n8868_o = n8774_o;
      6'b001000: n8868_o = n8583_o;
      6'b000100: n8868_o = ip;
      6'b000010: n8868_o = ip;
      6'b000001: n8868_o = ip;
      default: n8868_o = ip;
    endcase
  assign n8869_o = n8585_o[0];
  assign n8870_o = n8798_o[0];
  assign n8871_o = psw[1];
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8872_o = n8871_o;
      6'b010000: n8872_o = n8870_o;
      6'b001000: n8872_o = n8869_o;
      6'b000100: n8872_o = n8871_o;
      6'b000010: n8872_o = n8871_o;
      6'b000001: n8872_o = n8871_o;
      default: n8872_o = n8871_o;
    endcase
  assign n8873_o = n8585_o[1];
  assign n8874_o = n8798_o[1];
  assign n8875_o = psw[2];
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8876_o = n8822_o;
      6'b010000: n8876_o = n8874_o;
      6'b001000: n8876_o = n8873_o;
      6'b000100: n8876_o = new_ov_i;
      6'b000010: n8876_o = n8875_o;
      6'b000001: n8876_o = n8875_o;
      default: n8876_o = n8875_o;
    endcase
  assign n8877_o = n8585_o[4:2];
  assign n8878_o = n8798_o[4:2];
  assign n8879_o = psw[5:3];
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8880_o = n8879_o;
      6'b010000: n8880_o = n8878_o;
      6'b001000: n8880_o = n8877_o;
      6'b000100: n8880_o = n8879_o;
      6'b000010: n8880_o = n8879_o;
      6'b000001: n8880_o = n8879_o;
      default: n8880_o = n8879_o;
    endcase
  assign n8881_o = n8585_o[5];
  assign n8882_o = n8798_o[5];
  assign n8883_o = psw[6];
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8884_o = n8883_o;
      6'b010000: n8884_o = n8882_o;
      6'b001000: n8884_o = n8881_o;
      6'b000100: n8884_o = n8352_o;
      6'b000010: n8884_o = n8883_o;
      6'b000001: n8884_o = n8883_o;
      default: n8884_o = n8883_o;
    endcase
  assign n8885_o = n8585_o[6];
  assign n8886_o = psw[7];
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8887_o = n8824_o;
      6'b010000: n8887_o = n8800_o;
      6'b001000: n8887_o = n8885_o;
      6'b000100: n8887_o = n8351_o;
      6'b000010: n8887_o = n8886_o;
      6'b000001: n8887_o = n8886_o;
      default: n8887_o = n8886_o;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8888_o = n8825_o;
      6'b010000: n8888_o = n8778_o;
      6'b001000: n8888_o = n8586_o;
      6'b000100: n8888_o = s_data;
      6'b000010: n8888_o = s_data;
      6'b000001: n8888_o = acc;
      default: n8888_o = acc;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8889_o = n8826_o;
      6'b010000: n8889_o = n8779_o;
      6'b001000: n8889_o = n8587_o;
      6'b000100: n8889_o = b;
      6'b000010: n8889_o = b;
      6'b000001: n8889_o = b;
      default: n8889_o = b;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8890_o = tsel;
      6'b010000: n8890_o = tsel;
      6'b001000: n8890_o = n8588_o;
      6'b000100: n8890_o = tsel;
      6'b000010: n8890_o = tsel;
      6'b000001: n8890_o = tsel;
      default: n8890_o = tsel;
    endcase
  /* control_mem_rtl.vhd:971:9  */
  always @*
    case (n8829_o)
      6'b100000: n8891_o = ssel;
      6'b010000: n8891_o = ssel;
      6'b001000: n8891_o = n8589_o;
      6'b000100: n8891_o = ssel;
      6'b000010: n8891_o = ssel;
      6'b000001: n8891_o = ssel;
      default: n8891_o = ssel;
    endcase
  assign n8920_o = {n8887_o, n8884_o, n8880_o, n8876_o, n8872_o, s_p};
  /* control_mem_rtl.vhd:898:5  */
  assign n8928_o = reset ? 1'b0 : 1'b1;
  assign n8933_o = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
  /* control_mem_rtl.vhd:768:7  */
  assign n8996_o = cen ? n8129_o : s_help;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n8997_q <= 8'b00000000;
    else
      n8997_q <= n8996_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n8998_o = cen ? n8142_o : s_help16;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n8999_q <= 16'b0000000000000000;
    else
      n8999_q <= n8998_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9000_o = cen ? n8149_o : s_helpb;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9001_q <= 1'b0;
    else
      n9001_q <= n9000_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9002_o = cen & n8099_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9003_o = n9002_o ? rom_data_i : s_ir;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9004_q <= 8'b00000000;
    else
      n9004_q <= n9003_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9005_o = cen ? n8836_o : gprbit;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9006_q <= n8933_o;
    else
      n9006_q <= n9005_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9007_o = cen ? n8837_o : s_r0_b0;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9008_q <= 8'b00000000;
    else
      n9008_q <= n9007_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9009_o = cen ? n8838_o : s_r1_b0;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9010_q <= 8'b00000000;
    else
      n9010_q <= n9009_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9011_o = cen ? n8839_o : s_r0_b1;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9012_q <= 8'b00000000;
    else
      n9012_q <= n9011_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9013_o = cen ? n8840_o : s_r1_b1;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9014_q <= 8'b00000000;
    else
      n9014_q <= n9013_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9015_o = cen ? n8841_o : s_r0_b2;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9016_q <= 8'b00000000;
    else
      n9016_q <= n9015_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9017_o = cen ? n8842_o : s_r1_b2;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9018_q <= 8'b00000000;
    else
      n9018_q <= n9017_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9019_o = cen ? n8843_o : s_r0_b3;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9020_q <= 8'b00000000;
    else
      n9020_q <= n9019_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9021_o = cen ? n8844_o : s_r1_b3;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9022_q <= 8'b00000000;
    else
      n9022_q <= n9021_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9023_o = cen ? s_nextstate : state;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9024_q <= 3'b000;
    else
      n9024_q <= n9023_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9025_o = cen & ext0isr_en_i;
  /* control_mem_rtl.vhd:768:7  */
  assign n9026_o = n9025_o ? ext0isr_d_i : s_ext0isr_d;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9027_q <= 1'b0;
    else
      n9027_q <= n9026_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9028_o = cen & ext0isrh_en_i;
  /* control_mem_rtl.vhd:768:7  */
  assign n9029_o = n9028_o ? ext0isrh_d_i : s_ext0isrh_d;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9030_q <= 1'b0;
    else
      n9030_q <= n9029_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9031_o = cen & ext1isr_en_i;
  /* control_mem_rtl.vhd:768:7  */
  assign n9032_o = n9031_o ? ext1isr_d_i : s_ext1isr_d;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9033_q <= 1'b0;
    else
      n9033_q <= n9032_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9034_o = cen & ext1isrh_en_i;
  /* control_mem_rtl.vhd:768:7  */
  assign n9035_o = n9034_o ? ext1isrh_d_i : s_ext1isrh_d;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9036_q <= 1'b0;
    else
      n9036_q <= n9035_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9037_o = cen & s_intpre2_en;
  /* control_mem_rtl.vhd:768:7  */
  assign n9038_o = n9037_o ? s_intpre2_d : s_intpre2;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9039_q <= 1'b0;
    else
      n9039_q <= n9038_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9040_o = cen & s_inthigh_en;
  /* control_mem_rtl.vhd:768:7  */
  assign n9041_o = n9040_o ? s_inthigh_d : s_inthigh;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9042_q <= 1'b0;
    else
      n9042_q <= n9041_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9043_o = cen & s_intlow_en;
  /* control_mem_rtl.vhd:768:7  */
  assign n9044_o = n9043_o ? s_intlow_d : s_intlow;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9045_q <= 1'b0;
    else
      n9045_q <= n9044_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9046_o = cen ? s_intblock : s_intblock_o;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9047_q <= 1'b0;
    else
      n9047_q <= n9046_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9048_o = cen ? n8845_o : s_smodreg;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9049_q <= 1'b0;
    else
      n9049_q <= n9048_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9050_o = cen ? n8846_o : s_reload;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9051_q <= 8'b00000000;
    else
      n9051_q <= n9050_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9052_o = cen ? n8847_o : s_wt;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9053_q <= 2'b00;
    else
      n9053_q <= n9052_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9054_o = cen ? int0_i : s_int0_h1;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9055_q <= 1'b1;
    else
      n9055_q <= n9054_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9056_o = cen ? s_int0_h1 : s_int0_h2;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9057_q <= 1'b1;
    else
      n9057_q <= n9056_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9058_o = cen ? s_int0_h2 : s_int0_h3;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9059_q <= 1'b1;
    else
      n9059_q <= n9058_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9060_o = cen ? int1_i : s_int1_h1;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9061_q <= 1'b1;
    else
      n9061_q <= n9060_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9062_o = cen ? s_int1_h1 : s_int1_h2;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9063_q <= 1'b1;
    else
      n9063_q <= n9062_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9064_o = cen ? s_int1_h2 : s_int1_h3;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9065_q <= 1'b1;
    else
      n9065_q <= n9064_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9066_o = cen ? all_tf0_i : s_tf0_h1;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9067_q <= 1'b0;
    else
      n9067_q <= n9066_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9068_o = cen ? s_tf0_h1 : s_tf0_h2;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9069_q <= 1'b0;
    else
      n9069_q <= n9068_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9070_o = cen ? all_tf1_i : s_tf1_h1;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9071_q <= 1'b0;
    else
      n9071_q <= n9070_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9072_o = cen ? s_tf1_h1 : s_tf1_h2;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9073_q <= 1'b0;
    else
      n9073_q <= n9072_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9074_o = cen ? n7767_o : s_ri_h1;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9075_q <= 1'b0;
    else
      n9075_q <= n9074_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9076_o = cen ? s_ri_h1 : s_ri_h2;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9077_q <= 1'b0;
    else
      n9077_q <= n9076_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9078_o = cen ? n7768_o : s_ti_h1;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9079_q <= 1'b0;
    else
      n9079_q <= n9078_o;
  /* control_mem_rtl.vhd:554:5  */
  assign n9080_o = cen ? s_ti_h1 : s_ti_h2;
  /* control_mem_rtl.vhd:554:5  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9081_q <= 1'b0;
    else
      n9081_q <= n9080_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9084_o = cen ? p0_i : s_p0;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9085_q <= 8'b11111111;
    else
      n9085_q <= n9084_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9086_o = cen ? p1_i : s_p1;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9087_q <= 8'b11111111;
    else
      n9087_q <= n9086_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9088_o = cen ? p2_i : s_p2;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9089_q <= 8'b11111111;
    else
      n9089_q <= n9088_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9090_o = cen ? p3_i : s_p3;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9091_q <= 8'b11111111;
    else
      n9091_q <= n9090_o;
  /* control_mem_rtl.vhd:768:7  */
  assign n9092_o = cen ? pc_comb : pc;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9093_q <= 16'b0000000000000000;
    else
      n9093_q <= n9092_o;
  /* control_mem_rtl.vhd:748:5  */
  assign n9094_o = {n8271_o, n8261_o, n8251_o};
  assign n9095_o = {n7949_o, n7935_o};
  /* control_mem_rtl.vhd:768:7  */
  assign n9096_o = cen ? s_adr : s_preadr;
  /* control_mem_rtl.vhd:768:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9097_q <= 8'b00000000;
    else
      n9097_q <= n9096_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9098_o = cen ? n8848_o : p0;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9099_q <= 8'b11111111;
    else
      n9099_q <= n9098_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9100_o = cen ? n8849_o : sp;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9101_q <= 8'b00000111;
    else
      n9101_q <= n9100_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9102_o = cen ? n8850_o : dpl;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9103_q <= 8'b00000000;
    else
      n9103_q <= n9102_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9104_o = cen ? n8851_o : dph;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9105_q <= 8'b00000000;
    else
      n9105_q <= n9104_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9106_o = cen ? n8852_o : pcon;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9107_q <= 4'b0000;
    else
      n9107_q <= n9106_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9108_o = cen ? n8858_o : tcon;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9109_q <= 8'b00000000;
    else
      n9109_q <= n9108_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9110_o = cen ? n8859_o : tmod;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9111_q <= 8'b00000000;
    else
      n9111_q <= n9110_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9112_o = cen ? n8860_o : p1;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9113_q <= 8'b11111111;
    else
      n9113_q <= n9112_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9114_o = cen ? n8863_o : scon;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9115_q <= 8'b00000000;
    else
      n9115_q <= n9114_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9116_o = cen ? n8864_o : sbuf;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9117_q <= 8'b00000000;
    else
      n9117_q <= n9116_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9118_o = cen ? n8865_o : p2;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9119_q <= 8'b11111111;
    else
      n9119_q <= n9118_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9120_o = cen ? n8866_o : ie;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9121_q <= 8'b00000000;
    else
      n9121_q <= n9120_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9122_o = cen ? n8867_o : p3;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9123_q <= 8'b11111111;
    else
      n9123_q <= n9122_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9124_o = cen ? n8868_o : ip;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9125_q <= 8'b00000000;
    else
      n9125_q <= n9124_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9126_o = cen ? n8920_o : psw;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9127_q <= 8'b00000000;
    else
      n9127_q <= n9126_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9128_o = cen ? n8888_o : acc;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9129_q <= 8'b00000000;
    else
      n9129_q <= n9128_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9130_o = cen ? n8889_o : b;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9131_q <= 8'b00000000;
    else
      n9131_q <= n9130_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9132_o = cen ? n8890_o : tsel;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9133_q <= 8'b00000000;
    else
      n9133_q <= n9132_o;
  /* control_mem_rtl.vhd:951:7  */
  assign n9134_o = cen ? n8891_o : ssel;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9135_q <= 8'b00000000;
    else
      n9135_q <= n9134_o;
  /* control_mem_rtl.vhd:898:5  */
  assign n9136_o = {n7285_o, n7287_o};
  /* control_mem_rtl.vhd:951:7  */
  assign n9137_o = cen ? n8831_o : n9138_q;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9138_q <= 1'b0;
    else
      n9138_q <= n9137_o;
  /* control_mem_rtl.vhd:898:5  */
  assign n9139_o = {n7308_o, n7309_o, n7310_o, n7311_o, n7312_o, n7313_o};
  /* control_mem_rtl.vhd:951:7  */
  assign n9140_o = cen ? n8834_o : n9141_q;
  /* control_mem_rtl.vhd:951:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n9141_q <= 1'b0;
    else
      n9141_q <= n9140_o;
  /* control_mem_rtl.vhd:898:5  */
  assign n9142_o = {n8050_o, n8048_o};
  /* control_mem_.vhd:177:9  */
  assign n9144_o = gprbit[7:0];
  /* control_mem_.vhd:176:9  */
  assign n9145_o = gprbit[15:8];
  /* control_mem_.vhd:175:9  */
  assign n9146_o = gprbit[23:16];
  /* control_mem_.vhd:174:9  */
  assign n9147_o = gprbit[31:24];
  /* control_mem_.vhd:173:9  */
  assign n9148_o = gprbit[39:32];
  /* control_mem_.vhd:172:9  */
  assign n9149_o = gprbit[47:40];
  /* control_mem_.vhd:171:9  */
  assign n9150_o = gprbit[55:48];
  /* control_mem_.vhd:170:9  */
  assign n9151_o = gprbit[63:56];
  /* control_mem_.vhd:169:9  */
  assign n9152_o = gprbit[71:64];
  /* control_mem_.vhd:168:9  */
  assign n9153_o = gprbit[79:72];
  /* control_mem_.vhd:167:9  */
  assign n9154_o = gprbit[87:80];
  /* control_mem_.vhd:166:9  */
  assign n9155_o = gprbit[95:88];
  /* control_mem_.vhd:165:9  */
  assign n9156_o = gprbit[103:96];
  /* control_mem_.vhd:164:9  */
  assign n9157_o = gprbit[111:104];
  /* control_mem_.vhd:163:9  */
  assign n9158_o = gprbit[119:112];
  /* control_mem_.vhd:162:9  */
  assign n9159_o = gprbit[127:120];
  /* control_mem_rtl.vhd:443:33  */
  assign n9160_o = n7635_o[1:0];
  /* control_mem_rtl.vhd:443:33  */
  always @*
    case (n9160_o)
      2'b00: n9161_o = n9144_o;
      2'b01: n9161_o = n9145_o;
      2'b10: n9161_o = n9146_o;
      2'b11: n9161_o = n9147_o;
    endcase
  /* control_mem_rtl.vhd:443:33  */
  assign n9162_o = n7635_o[1:0];
  /* control_mem_rtl.vhd:443:33  */
  always @*
    case (n9162_o)
      2'b00: n9163_o = n9148_o;
      2'b01: n9163_o = n9149_o;
      2'b10: n9163_o = n9150_o;
      2'b11: n9163_o = n9151_o;
    endcase
  /* control_mem_rtl.vhd:443:33  */
  assign n9164_o = n7635_o[1:0];
  /* control_mem_rtl.vhd:443:33  */
  always @*
    case (n9164_o)
      2'b00: n9165_o = n9152_o;
      2'b01: n9165_o = n9153_o;
      2'b10: n9165_o = n9154_o;
      2'b11: n9165_o = n9155_o;
    endcase
  /* control_mem_rtl.vhd:443:33  */
  assign n9166_o = n7635_o[1:0];
  /* control_mem_rtl.vhd:443:33  */
  always @*
    case (n9166_o)
      2'b00: n9167_o = n9156_o;
      2'b01: n9167_o = n9157_o;
      2'b10: n9167_o = n9158_o;
      2'b11: n9167_o = n9159_o;
    endcase
  /* control_mem_rtl.vhd:443:33  */
  assign n9168_o = n7635_o[3:2];
  /* control_mem_rtl.vhd:443:33  */
  always @*
    case (n9168_o)
      2'b00: n9169_o = n9161_o;
      2'b01: n9169_o = n9163_o;
      2'b10: n9169_o = n9165_o;
      2'b11: n9169_o = n9167_o;
    endcase
  /* control_mem_rtl.vhd:443:33  */
  assign n9170_o = s_p0[0];
  /* control_mem_rtl.vhd:443:34  */
  assign n9171_o = s_p0[1];
  /* control_mem_.vhd:132:9  */
  assign n9172_o = s_p0[2];
  /* control_mem_.vhd:130:9  */
  assign n9173_o = s_p0[3];
  /* control_mem_.vhd:121:9  */
  assign n9174_o = s_p0[4];
  /* control_mem_.vhd:119:9  */
  assign n9175_o = s_p0[5];
  /* control_mem_.vhd:117:9  */
  assign n9176_o = s_p0[6];
  /* control_mem_.vhd:115:9  */
  assign n9177_o = s_p0[7];
  /* control_mem_rtl.vhd:468:42  */
  assign n9178_o = n7668_o[1:0];
  /* control_mem_rtl.vhd:468:42  */
  always @*
    case (n9178_o)
      2'b00: n9179_o = n9170_o;
      2'b01: n9179_o = n9171_o;
      2'b10: n9179_o = n9172_o;
      2'b11: n9179_o = n9173_o;
    endcase
  /* control_mem_rtl.vhd:468:42  */
  assign n9180_o = n7668_o[1:0];
  /* control_mem_rtl.vhd:468:42  */
  always @*
    case (n9180_o)
      2'b00: n9181_o = n9174_o;
      2'b01: n9181_o = n9175_o;
      2'b10: n9181_o = n9176_o;
      2'b11: n9181_o = n9177_o;
    endcase
  /* control_mem_rtl.vhd:468:42  */
  assign n9182_o = n7668_o[2];
  /* control_mem_rtl.vhd:468:42  */
  assign n9183_o = n9182_o ? n9181_o : n9179_o;
  /* control_mem_rtl.vhd:468:42  */
  assign n9184_o = tcon[0];
  /* control_mem_rtl.vhd:468:43  */
  assign n9185_o = tcon[1];
  /* control_mem_.vhd:89:9  */
  assign n9186_o = tcon[2];
  /* control_mem_.vhd:88:9  */
  assign n9187_o = tcon[3];
  /* control_mem_.vhd:86:9  */
  assign n9188_o = tcon[4];
  /* control_mem_.vhd:85:9  */
  assign n9189_o = tcon[5];
  /* control_mem_.vhd:84:9  */
  assign n9190_o = tcon[6];
  /* control_mem_.vhd:80:9  */
  assign n9191_o = tcon[7];
  /* control_mem_rtl.vhd:470:37  */
  assign n9192_o = n7674_o[1:0];
  /* control_mem_rtl.vhd:470:37  */
  always @*
    case (n9192_o)
      2'b00: n9193_o = n9184_o;
      2'b01: n9193_o = n9185_o;
      2'b10: n9193_o = n9186_o;
      2'b11: n9193_o = n9187_o;
    endcase
  /* control_mem_rtl.vhd:470:37  */
  assign n9194_o = n7674_o[1:0];
  /* control_mem_rtl.vhd:470:37  */
  always @*
    case (n9194_o)
      2'b00: n9195_o = n9188_o;
      2'b01: n9195_o = n9189_o;
      2'b10: n9195_o = n9190_o;
      2'b11: n9195_o = n9191_o;
    endcase
  /* control_mem_rtl.vhd:470:37  */
  assign n9196_o = n7674_o[2];
  /* control_mem_rtl.vhd:470:37  */
  assign n9197_o = n9196_o ? n9195_o : n9193_o;
  /* control_mem_rtl.vhd:470:37  */
  assign n9198_o = s_p1[0];
  /* control_mem_rtl.vhd:470:38  */
  assign n9199_o = s_p1[1];
  assign n9200_o = s_p1[2];
  /* control_mem_rtl.vhd:1124:24  */
  assign n9201_o = s_p1[3];
  /* control_mem_rtl.vhd:1123:24  */
  assign n9202_o = s_p1[4];
  /* control_mem_rtl.vhd:1119:23  */
  assign n9203_o = s_p1[5];
  /* control_mem_rtl.vhd:1117:25  */
  assign n9204_o = s_p1[6];
  /* control_mem_rtl.vhd:1103:24  */
  assign n9205_o = s_p1[7];
  /* control_mem_rtl.vhd:471:42  */
  assign n9206_o = n7680_o[1:0];
  /* control_mem_rtl.vhd:471:42  */
  always @*
    case (n9206_o)
      2'b00: n9207_o = n9198_o;
      2'b01: n9207_o = n9199_o;
      2'b10: n9207_o = n9200_o;
      2'b11: n9207_o = n9201_o;
    endcase
  /* control_mem_rtl.vhd:471:42  */
  assign n9208_o = n7680_o[1:0];
  /* control_mem_rtl.vhd:471:42  */
  always @*
    case (n9208_o)
      2'b00: n9209_o = n9202_o;
      2'b01: n9209_o = n9203_o;
      2'b10: n9209_o = n9204_o;
      2'b11: n9209_o = n9205_o;
    endcase
  /* control_mem_rtl.vhd:471:42  */
  assign n9210_o = n7680_o[2];
  /* control_mem_rtl.vhd:471:42  */
  assign n9211_o = n9210_o ? n9209_o : n9207_o;
  /* control_mem_rtl.vhd:471:42  */
  assign n9212_o = scon[0];
  /* control_mem_rtl.vhd:471:43  */
  assign n9213_o = scon[1];
  /* control_mem_rtl.vhd:1089:24  */
  assign n9214_o = scon[2];
  /* control_mem_rtl.vhd:1059:22  */
  assign n9215_o = scon[3];
  assign n9216_o = scon[4];
  assign n9217_o = scon[5];
  assign n9218_o = scon[6];
  assign n9219_o = scon[7];
  /* control_mem_rtl.vhd:476:39  */
  assign n9220_o = n7690_o[1:0];
  /* control_mem_rtl.vhd:476:39  */
  always @*
    case (n9220_o)
      2'b00: n9221_o = n9212_o;
      2'b01: n9221_o = n9213_o;
      2'b10: n9221_o = n9214_o;
      2'b11: n9221_o = n9215_o;
    endcase
  /* control_mem_rtl.vhd:476:39  */
  assign n9222_o = n7690_o[1:0];
  /* control_mem_rtl.vhd:476:39  */
  always @*
    case (n9222_o)
      2'b00: n9223_o = n9216_o;
      2'b01: n9223_o = n9217_o;
      2'b10: n9223_o = n9218_o;
      2'b11: n9223_o = n9219_o;
    endcase
  /* control_mem_rtl.vhd:476:39  */
  assign n9224_o = n7690_o[2];
  /* control_mem_rtl.vhd:476:39  */
  assign n9225_o = n9224_o ? n9223_o : n9221_o;
  /* control_mem_rtl.vhd:476:39  */
  assign n9226_o = s_p2[0];
  /* control_mem_rtl.vhd:476:40  */
  assign n9227_o = s_p2[1];
  /* control_mem_rtl.vhd:856:3  */
  assign n9228_o = s_p2[2];
  /* control_mem_rtl.vhd:858:12  */
  assign n9229_o = s_p2[3];
  assign n9230_o = s_p2[4];
  assign n9231_o = s_p2[5];
  /* control_mem_rtl.vhd:768:7  */
  assign n9232_o = s_p2[6];
  /* control_mem_rtl.vhd:768:7  */
  assign n9233_o = s_p2[7];
  /* control_mem_rtl.vhd:478:42  */
  assign n9234_o = n7697_o[1:0];
  /* control_mem_rtl.vhd:478:42  */
  always @*
    case (n9234_o)
      2'b00: n9235_o = n9226_o;
      2'b01: n9235_o = n9227_o;
      2'b10: n9235_o = n9228_o;
      2'b11: n9235_o = n9229_o;
    endcase
  /* control_mem_rtl.vhd:478:42  */
  assign n9236_o = n7697_o[1:0];
  /* control_mem_rtl.vhd:478:42  */
  always @*
    case (n9236_o)
      2'b00: n9237_o = n9230_o;
      2'b01: n9237_o = n9231_o;
      2'b10: n9237_o = n9232_o;
      2'b11: n9237_o = n9233_o;
    endcase
  /* control_mem_rtl.vhd:478:42  */
  assign n9238_o = n7697_o[2];
  /* control_mem_rtl.vhd:478:42  */
  assign n9239_o = n9238_o ? n9237_o : n9235_o;
  /* control_mem_rtl.vhd:478:42  */
  assign n9240_o = ie[0];
  /* control_mem_rtl.vhd:478:43  */
  assign n9241_o = ie[1];
  assign n9242_o = ie[2];
  /* control_mem_rtl.vhd:768:27  */
  assign n9243_o = ie[3];
  /* control_mem_rtl.vhd:746:3  */
  assign n9244_o = ie[4];
  assign n9245_o = ie[5];
  assign n9246_o = ie[6];
  /* control_mem_rtl.vhd:630:3  */
  assign n9247_o = ie[7];
  /* control_mem_rtl.vhd:479:40  */
  assign n9248_o = n7703_o[1:0];
  /* control_mem_rtl.vhd:479:40  */
  always @*
    case (n9248_o)
      2'b00: n9249_o = n9240_o;
      2'b01: n9249_o = n9241_o;
      2'b10: n9249_o = n9242_o;
      2'b11: n9249_o = n9243_o;
    endcase
  /* control_mem_rtl.vhd:479:40  */
  assign n9250_o = n7703_o[1:0];
  /* control_mem_rtl.vhd:479:40  */
  always @*
    case (n9250_o)
      2'b00: n9251_o = n9244_o;
      2'b01: n9251_o = n9245_o;
      2'b10: n9251_o = n9246_o;
      2'b11: n9251_o = n9247_o;
    endcase
  /* control_mem_rtl.vhd:479:40  */
  assign n9252_o = n7703_o[2];
  /* control_mem_rtl.vhd:479:40  */
  assign n9253_o = n9252_o ? n9251_o : n9249_o;
  /* control_mem_rtl.vhd:479:40  */
  assign n9254_o = s_p3[0];
  /* control_mem_rtl.vhd:479:41  */
  assign n9255_o = s_p3[1];
  /* control_mem_rtl.vhd:489:28  */
  assign n9256_o = s_p3[2];
  /* control_mem_rtl.vhd:488:34  */
  assign n9257_o = s_p3[3];
  /* control_mem_rtl.vhd:484:40  */
  assign n9258_o = s_p3[4];
  /* control_mem_rtl.vhd:483:42  */
  assign n9259_o = s_p3[5];
  /* control_mem_rtl.vhd:482:42  */
  assign n9260_o = s_p3[6];
  /* control_mem_rtl.vhd:481:41  */
  assign n9261_o = s_p3[7];
  /* control_mem_rtl.vhd:480:42  */
  assign n9262_o = n7709_o[1:0];
  /* control_mem_rtl.vhd:480:42  */
  always @*
    case (n9262_o)
      2'b00: n9263_o = n9254_o;
      2'b01: n9263_o = n9255_o;
      2'b10: n9263_o = n9256_o;
      2'b11: n9263_o = n9257_o;
    endcase
  /* control_mem_rtl.vhd:480:42  */
  assign n9264_o = n7709_o[1:0];
  /* control_mem_rtl.vhd:480:42  */
  always @*
    case (n9264_o)
      2'b00: n9265_o = n9258_o;
      2'b01: n9265_o = n9259_o;
      2'b10: n9265_o = n9260_o;
      2'b11: n9265_o = n9261_o;
    endcase
  /* control_mem_rtl.vhd:480:42  */
  assign n9266_o = n7709_o[2];
  /* control_mem_rtl.vhd:480:42  */
  assign n9267_o = n9266_o ? n9265_o : n9263_o;
  /* control_mem_rtl.vhd:480:42  */
  assign n9268_o = ip[0];
  /* control_mem_rtl.vhd:480:43  */
  assign n9269_o = ip[1];
  /* control_mem_rtl.vhd:468:43  */
  assign n9270_o = ip[2];
  /* control_mem_rtl.vhd:443:34  */
  assign n9271_o = ip[3];
  /* control_mem_rtl.vhd:396:3  */
  assign n9272_o = ip[4];
  assign n9273_o = ip[5];
  /* control_mem_rtl.vhd:364:5  */
  assign n9274_o = ip[6];
  assign n9275_o = ip[7];
  /* control_mem_rtl.vhd:481:40  */
  assign n9276_o = n7715_o[1:0];
  /* control_mem_rtl.vhd:481:40  */
  always @*
    case (n9276_o)
      2'b00: n9277_o = n9268_o;
      2'b01: n9277_o = n9269_o;
      2'b10: n9277_o = n9270_o;
      2'b11: n9277_o = n9271_o;
    endcase
  /* control_mem_rtl.vhd:481:40  */
  assign n9278_o = n7715_o[1:0];
  /* control_mem_rtl.vhd:481:40  */
  always @*
    case (n9278_o)
      2'b00: n9279_o = n9272_o;
      2'b01: n9279_o = n9273_o;
      2'b10: n9279_o = n9274_o;
      2'b11: n9279_o = n9275_o;
    endcase
  /* control_mem_rtl.vhd:481:40  */
  assign n9280_o = n7715_o[2];
  /* control_mem_rtl.vhd:481:40  */
  assign n9281_o = n9280_o ? n9279_o : n9277_o;
  /* control_mem_rtl.vhd:481:40  */
  assign n9282_o = psw[0];
  /* control_mem_rtl.vhd:481:41  */
  assign n9283_o = psw[1];
  assign n9284_o = psw[2];
  /* control_mem_rtl.vhd:278:32  */
  assign n9285_o = psw[3];
  /* control_mem_rtl.vhd:278:42  */
  assign n9286_o = psw[4];
  /* control_mem_rtl.vhd:278:42  */
  assign n9287_o = psw[5];
  /* control_mem_rtl.vhd:278:42  */
  assign n9288_o = psw[6];
  /* control_mem_rtl.vhd:278:13  */
  assign n9289_o = psw[7];
  /* control_mem_rtl.vhd:482:41  */
  assign n9290_o = n7721_o[1:0];
  /* control_mem_rtl.vhd:482:41  */
  always @*
    case (n9290_o)
      2'b00: n9291_o = n9282_o;
      2'b01: n9291_o = n9283_o;
      2'b10: n9291_o = n9284_o;
      2'b11: n9291_o = n9285_o;
    endcase
  /* control_mem_rtl.vhd:482:41  */
  assign n9292_o = n7721_o[1:0];
  /* control_mem_rtl.vhd:482:41  */
  always @*
    case (n9292_o)
      2'b00: n9293_o = n9286_o;
      2'b01: n9293_o = n9287_o;
      2'b10: n9293_o = n9288_o;
      2'b11: n9293_o = n9289_o;
    endcase
  /* control_mem_rtl.vhd:482:41  */
  assign n9294_o = n7721_o[2];
  /* control_mem_rtl.vhd:482:41  */
  assign n9295_o = n9294_o ? n9293_o : n9291_o;
  /* control_mem_rtl.vhd:482:41  */
  assign n9296_o = acc[0];
  /* control_mem_rtl.vhd:482:42  */
  assign n9297_o = acc[1];
  assign n9298_o = acc[2];
  assign n9299_o = acc[3];
  assign n9300_o = acc[4];
  assign n9301_o = acc[5];
  assign n9302_o = acc[6];
  assign n9303_o = acc[7];
  /* control_mem_rtl.vhd:483:41  */
  assign n9304_o = n7727_o[1:0];
  /* control_mem_rtl.vhd:483:41  */
  always @*
    case (n9304_o)
      2'b00: n9305_o = n9296_o;
      2'b01: n9305_o = n9297_o;
      2'b10: n9305_o = n9298_o;
      2'b11: n9305_o = n9299_o;
    endcase
  /* control_mem_rtl.vhd:483:41  */
  assign n9306_o = n7727_o[1:0];
  /* control_mem_rtl.vhd:483:41  */
  always @*
    case (n9306_o)
      2'b00: n9307_o = n9300_o;
      2'b01: n9307_o = n9301_o;
      2'b10: n9307_o = n9302_o;
      2'b11: n9307_o = n9303_o;
    endcase
  /* control_mem_rtl.vhd:483:41  */
  assign n9308_o = n7727_o[2];
  /* control_mem_rtl.vhd:483:41  */
  assign n9309_o = n9308_o ? n9307_o : n9305_o;
  /* control_mem_rtl.vhd:483:41  */
  assign n9310_o = b[0];
  /* control_mem_rtl.vhd:483:42  */
  assign n9311_o = b[1];
  assign n9312_o = b[2];
  assign n9313_o = b[3];
  assign n9314_o = b[4];
  assign n9315_o = b[5];
  assign n9316_o = b[6];
  assign n9317_o = b[7];
  /* control_mem_rtl.vhd:484:39  */
  assign n9318_o = n7733_o[1:0];
  /* control_mem_rtl.vhd:484:39  */
  always @*
    case (n9318_o)
      2'b00: n9319_o = n9310_o;
      2'b01: n9319_o = n9311_o;
      2'b10: n9319_o = n9312_o;
      2'b11: n9319_o = n9313_o;
    endcase
  /* control_mem_rtl.vhd:484:39  */
  assign n9320_o = n7733_o[1:0];
  /* control_mem_rtl.vhd:484:39  */
  always @*
    case (n9320_o)
      2'b00: n9321_o = n9314_o;
      2'b01: n9321_o = n9315_o;
      2'b10: n9321_o = n9316_o;
      2'b11: n9321_o = n9317_o;
    endcase
  /* control_mem_rtl.vhd:484:39  */
  assign n9322_o = n7733_o[2];
  /* control_mem_rtl.vhd:484:39  */
  assign n9323_o = n9322_o ? n9321_o : n9319_o;
  /* control_mem_rtl.vhd:484:39  */
  assign n9324_o = gprbit[0];
  /* control_mem_rtl.vhd:484:40  */
  assign n9325_o = gprbit[1];
  assign n9326_o = gprbit[2];
  assign n9327_o = gprbit[3];
  assign n9328_o = gprbit[4];
  assign n9329_o = gprbit[5];
  assign n9330_o = gprbit[6];
  assign n9331_o = gprbit[7];
  assign n9332_o = gprbit[8];
  assign n9333_o = gprbit[9];
  assign n9334_o = gprbit[10];
  assign n9335_o = gprbit[11];
  assign n9336_o = gprbit[12];
  assign n9337_o = gprbit[13];
  assign n9338_o = gprbit[14];
  assign n9339_o = gprbit[15];
  assign n9340_o = gprbit[16];
  assign n9341_o = gprbit[17];
  assign n9342_o = gprbit[18];
  assign n9343_o = gprbit[19];
  assign n9344_o = gprbit[20];
  assign n9345_o = gprbit[21];
  assign n9346_o = gprbit[22];
  assign n9347_o = gprbit[23];
  assign n9348_o = gprbit[24];
  assign n9349_o = gprbit[25];
  assign n9350_o = gprbit[26];
  assign n9351_o = gprbit[27];
  assign n9352_o = gprbit[28];
  assign n9353_o = gprbit[29];
  assign n9354_o = gprbit[30];
  assign n9355_o = gprbit[31];
  assign n9356_o = gprbit[32];
  assign n9357_o = gprbit[33];
  assign n9358_o = gprbit[34];
  assign n9359_o = gprbit[35];
  assign n9360_o = gprbit[36];
  assign n9361_o = gprbit[37];
  assign n9362_o = gprbit[38];
  assign n9363_o = gprbit[39];
  assign n9364_o = gprbit[40];
  assign n9365_o = gprbit[41];
  assign n9366_o = gprbit[42];
  assign n9367_o = gprbit[43];
  assign n9368_o = gprbit[44];
  assign n9369_o = gprbit[45];
  assign n9370_o = gprbit[46];
  assign n9371_o = gprbit[47];
  assign n9372_o = gprbit[48];
  assign n9373_o = gprbit[49];
  assign n9374_o = gprbit[50];
  assign n9375_o = gprbit[51];
  assign n9376_o = gprbit[52];
  assign n9377_o = gprbit[53];
  assign n9378_o = gprbit[54];
  assign n9379_o = gprbit[55];
  assign n9380_o = gprbit[56];
  assign n9381_o = gprbit[57];
  assign n9382_o = gprbit[58];
  assign n9383_o = gprbit[59];
  assign n9384_o = gprbit[60];
  assign n9385_o = gprbit[61];
  assign n9386_o = gprbit[62];
  assign n9387_o = gprbit[63];
  assign n9388_o = gprbit[64];
  assign n9389_o = gprbit[65];
  assign n9390_o = gprbit[66];
  assign n9391_o = gprbit[67];
  assign n9392_o = gprbit[68];
  assign n9393_o = gprbit[69];
  assign n9394_o = gprbit[70];
  assign n9395_o = gprbit[71];
  assign n9396_o = gprbit[72];
  assign n9397_o = gprbit[73];
  assign n9398_o = gprbit[74];
  assign n9399_o = gprbit[75];
  assign n9400_o = gprbit[76];
  assign n9401_o = gprbit[77];
  assign n9402_o = gprbit[78];
  assign n9403_o = gprbit[79];
  assign n9404_o = gprbit[80];
  assign n9405_o = gprbit[81];
  assign n9406_o = gprbit[82];
  assign n9407_o = gprbit[83];
  assign n9408_o = gprbit[84];
  assign n9409_o = gprbit[85];
  assign n9410_o = gprbit[86];
  assign n9411_o = gprbit[87];
  assign n9412_o = gprbit[88];
  assign n9413_o = gprbit[89];
  assign n9414_o = gprbit[90];
  assign n9415_o = gprbit[91];
  assign n9416_o = gprbit[92];
  assign n9417_o = gprbit[93];
  assign n9418_o = gprbit[94];
  assign n9419_o = gprbit[95];
  assign n9420_o = gprbit[96];
  assign n9421_o = gprbit[97];
  assign n9422_o = gprbit[98];
  assign n9423_o = gprbit[99];
  assign n9424_o = gprbit[100];
  assign n9425_o = gprbit[101];
  assign n9426_o = gprbit[102];
  assign n9427_o = gprbit[103];
  assign n9428_o = gprbit[104];
  assign n9429_o = gprbit[105];
  assign n9430_o = gprbit[106];
  assign n9431_o = gprbit[107];
  assign n9432_o = gprbit[108];
  assign n9433_o = gprbit[109];
  assign n9434_o = gprbit[110];
  assign n9435_o = gprbit[111];
  assign n9436_o = gprbit[112];
  assign n9437_o = gprbit[113];
  assign n9438_o = gprbit[114];
  assign n9439_o = gprbit[115];
  assign n9440_o = gprbit[116];
  assign n9441_o = gprbit[117];
  assign n9442_o = gprbit[118];
  assign n9443_o = gprbit[119];
  assign n9444_o = gprbit[120];
  assign n9445_o = gprbit[121];
  assign n9446_o = gprbit[122];
  assign n9447_o = gprbit[123];
  assign n9448_o = gprbit[124];
  assign n9449_o = gprbit[125];
  assign n9450_o = gprbit[126];
  assign n9451_o = gprbit[127];
  /* control_mem_rtl.vhd:489:27  */
  assign n9452_o = {n7742_o, n7745_o};
  /* control_mem_rtl.vhd:489:27  */
  assign n9453_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9453_o)
      2'b00: n9454_o = n9324_o;
      2'b01: n9454_o = n9325_o;
      2'b10: n9454_o = n9326_o;
      2'b11: n9454_o = n9327_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9455_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9455_o)
      2'b00: n9456_o = n9328_o;
      2'b01: n9456_o = n9329_o;
      2'b10: n9456_o = n9330_o;
      2'b11: n9456_o = n9331_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9457_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9457_o)
      2'b00: n9458_o = n9332_o;
      2'b01: n9458_o = n9333_o;
      2'b10: n9458_o = n9334_o;
      2'b11: n9458_o = n9335_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9459_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9459_o)
      2'b00: n9460_o = n9336_o;
      2'b01: n9460_o = n9337_o;
      2'b10: n9460_o = n9338_o;
      2'b11: n9460_o = n9339_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9461_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9461_o)
      2'b00: n9462_o = n9340_o;
      2'b01: n9462_o = n9341_o;
      2'b10: n9462_o = n9342_o;
      2'b11: n9462_o = n9343_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9463_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9463_o)
      2'b00: n9464_o = n9344_o;
      2'b01: n9464_o = n9345_o;
      2'b10: n9464_o = n9346_o;
      2'b11: n9464_o = n9347_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9465_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9465_o)
      2'b00: n9466_o = n9348_o;
      2'b01: n9466_o = n9349_o;
      2'b10: n9466_o = n9350_o;
      2'b11: n9466_o = n9351_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9467_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9467_o)
      2'b00: n9468_o = n9352_o;
      2'b01: n9468_o = n9353_o;
      2'b10: n9468_o = n9354_o;
      2'b11: n9468_o = n9355_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9469_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9469_o)
      2'b00: n9470_o = n9356_o;
      2'b01: n9470_o = n9357_o;
      2'b10: n9470_o = n9358_o;
      2'b11: n9470_o = n9359_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9471_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9471_o)
      2'b00: n9472_o = n9360_o;
      2'b01: n9472_o = n9361_o;
      2'b10: n9472_o = n9362_o;
      2'b11: n9472_o = n9363_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9473_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9473_o)
      2'b00: n9474_o = n9364_o;
      2'b01: n9474_o = n9365_o;
      2'b10: n9474_o = n9366_o;
      2'b11: n9474_o = n9367_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9475_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9475_o)
      2'b00: n9476_o = n9368_o;
      2'b01: n9476_o = n9369_o;
      2'b10: n9476_o = n9370_o;
      2'b11: n9476_o = n9371_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9477_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9477_o)
      2'b00: n9478_o = n9372_o;
      2'b01: n9478_o = n9373_o;
      2'b10: n9478_o = n9374_o;
      2'b11: n9478_o = n9375_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9479_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9479_o)
      2'b00: n9480_o = n9376_o;
      2'b01: n9480_o = n9377_o;
      2'b10: n9480_o = n9378_o;
      2'b11: n9480_o = n9379_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9481_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9481_o)
      2'b00: n9482_o = n9380_o;
      2'b01: n9482_o = n9381_o;
      2'b10: n9482_o = n9382_o;
      2'b11: n9482_o = n9383_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9483_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9483_o)
      2'b00: n9484_o = n9384_o;
      2'b01: n9484_o = n9385_o;
      2'b10: n9484_o = n9386_o;
      2'b11: n9484_o = n9387_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9485_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9485_o)
      2'b00: n9486_o = n9388_o;
      2'b01: n9486_o = n9389_o;
      2'b10: n9486_o = n9390_o;
      2'b11: n9486_o = n9391_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9487_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9487_o)
      2'b00: n9488_o = n9392_o;
      2'b01: n9488_o = n9393_o;
      2'b10: n9488_o = n9394_o;
      2'b11: n9488_o = n9395_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9489_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9489_o)
      2'b00: n9490_o = n9396_o;
      2'b01: n9490_o = n9397_o;
      2'b10: n9490_o = n9398_o;
      2'b11: n9490_o = n9399_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9491_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9491_o)
      2'b00: n9492_o = n9400_o;
      2'b01: n9492_o = n9401_o;
      2'b10: n9492_o = n9402_o;
      2'b11: n9492_o = n9403_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9493_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9493_o)
      2'b00: n9494_o = n9404_o;
      2'b01: n9494_o = n9405_o;
      2'b10: n9494_o = n9406_o;
      2'b11: n9494_o = n9407_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9495_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9495_o)
      2'b00: n9496_o = n9408_o;
      2'b01: n9496_o = n9409_o;
      2'b10: n9496_o = n9410_o;
      2'b11: n9496_o = n9411_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9497_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9497_o)
      2'b00: n9498_o = n9412_o;
      2'b01: n9498_o = n9413_o;
      2'b10: n9498_o = n9414_o;
      2'b11: n9498_o = n9415_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9499_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9499_o)
      2'b00: n9500_o = n9416_o;
      2'b01: n9500_o = n9417_o;
      2'b10: n9500_o = n9418_o;
      2'b11: n9500_o = n9419_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9501_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9501_o)
      2'b00: n9502_o = n9420_o;
      2'b01: n9502_o = n9421_o;
      2'b10: n9502_o = n9422_o;
      2'b11: n9502_o = n9423_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9503_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9503_o)
      2'b00: n9504_o = n9424_o;
      2'b01: n9504_o = n9425_o;
      2'b10: n9504_o = n9426_o;
      2'b11: n9504_o = n9427_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9505_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9505_o)
      2'b00: n9506_o = n9428_o;
      2'b01: n9506_o = n9429_o;
      2'b10: n9506_o = n9430_o;
      2'b11: n9506_o = n9431_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9507_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9507_o)
      2'b00: n9508_o = n9432_o;
      2'b01: n9508_o = n9433_o;
      2'b10: n9508_o = n9434_o;
      2'b11: n9508_o = n9435_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9509_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9509_o)
      2'b00: n9510_o = n9436_o;
      2'b01: n9510_o = n9437_o;
      2'b10: n9510_o = n9438_o;
      2'b11: n9510_o = n9439_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9511_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9511_o)
      2'b00: n9512_o = n9440_o;
      2'b01: n9512_o = n9441_o;
      2'b10: n9512_o = n9442_o;
      2'b11: n9512_o = n9443_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9513_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9513_o)
      2'b00: n9514_o = n9444_o;
      2'b01: n9514_o = n9445_o;
      2'b10: n9514_o = n9446_o;
      2'b11: n9514_o = n9447_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9515_o = n9452_o[1:0];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9515_o)
      2'b00: n9516_o = n9448_o;
      2'b01: n9516_o = n9449_o;
      2'b10: n9516_o = n9450_o;
      2'b11: n9516_o = n9451_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9517_o = n9452_o[3:2];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9517_o)
      2'b00: n9518_o = n9454_o;
      2'b01: n9518_o = n9456_o;
      2'b10: n9518_o = n9458_o;
      2'b11: n9518_o = n9460_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9519_o = n9452_o[3:2];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9519_o)
      2'b00: n9520_o = n9462_o;
      2'b01: n9520_o = n9464_o;
      2'b10: n9520_o = n9466_o;
      2'b11: n9520_o = n9468_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9521_o = n9452_o[3:2];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9521_o)
      2'b00: n9522_o = n9470_o;
      2'b01: n9522_o = n9472_o;
      2'b10: n9522_o = n9474_o;
      2'b11: n9522_o = n9476_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9523_o = n9452_o[3:2];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9523_o)
      2'b00: n9524_o = n9478_o;
      2'b01: n9524_o = n9480_o;
      2'b10: n9524_o = n9482_o;
      2'b11: n9524_o = n9484_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9525_o = n9452_o[3:2];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9525_o)
      2'b00: n9526_o = n9486_o;
      2'b01: n9526_o = n9488_o;
      2'b10: n9526_o = n9490_o;
      2'b11: n9526_o = n9492_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9527_o = n9452_o[3:2];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9527_o)
      2'b00: n9528_o = n9494_o;
      2'b01: n9528_o = n9496_o;
      2'b10: n9528_o = n9498_o;
      2'b11: n9528_o = n9500_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9529_o = n9452_o[3:2];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9529_o)
      2'b00: n9530_o = n9502_o;
      2'b01: n9530_o = n9504_o;
      2'b10: n9530_o = n9506_o;
      2'b11: n9530_o = n9508_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9531_o = n9452_o[3:2];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9531_o)
      2'b00: n9532_o = n9510_o;
      2'b01: n9532_o = n9512_o;
      2'b10: n9532_o = n9514_o;
      2'b11: n9532_o = n9516_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9533_o = n9452_o[5:4];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9533_o)
      2'b00: n9534_o = n9518_o;
      2'b01: n9534_o = n9520_o;
      2'b10: n9534_o = n9522_o;
      2'b11: n9534_o = n9524_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9535_o = n9452_o[5:4];
  /* control_mem_rtl.vhd:489:27  */
  always @*
    case (n9535_o)
      2'b00: n9536_o = n9526_o;
      2'b01: n9536_o = n9528_o;
      2'b10: n9536_o = n9530_o;
      2'b11: n9536_o = n9532_o;
    endcase
  /* control_mem_rtl.vhd:489:27  */
  assign n9537_o = n9452_o[6];
  /* control_mem_rtl.vhd:489:27  */
  assign n9538_o = n9537_o ? n9536_o : n9534_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9539_o = n8483_o[3];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9540_o = ~n9539_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9541_o = n8483_o[2];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9542_o = ~n9541_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9543_o = n9540_o & n9542_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9544_o = n9540_o & n9541_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9545_o = n9539_o & n9542_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9546_o = n9539_o & n9541_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9547_o = n8483_o[1];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9548_o = ~n9547_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9549_o = n9543_o & n9548_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9550_o = n9543_o & n9547_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9551_o = n9544_o & n9548_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9552_o = n9544_o & n9547_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9553_o = n9545_o & n9548_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9554_o = n9545_o & n9547_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9555_o = n9546_o & n9548_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9556_o = n9546_o & n9547_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9557_o = n8483_o[0];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9558_o = ~n9557_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9559_o = n9549_o & n9558_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9560_o = n9549_o & n9557_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9561_o = n9550_o & n9558_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9562_o = n9550_o & n9557_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9563_o = n9551_o & n9558_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9564_o = n9551_o & n9557_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9565_o = n9552_o & n9558_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9566_o = n9552_o & n9557_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9567_o = n9553_o & n9558_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9568_o = n9553_o & n9557_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9569_o = n9554_o & n9558_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9570_o = n9554_o & n9557_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9571_o = n9555_o & n9558_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9572_o = n9555_o & n9557_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9573_o = n9556_o & n9558_o;
  /* control_mem_rtl.vhd:1059:15  */
  assign n9574_o = n9556_o & n9557_o;
  assign n9575_o = gprbit[7:0];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9576_o = n9559_o ? s_data : n9575_o;
  assign n9577_o = gprbit[15:8];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9578_o = n9560_o ? s_data : n9577_o;
  assign n9579_o = gprbit[23:16];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9580_o = n9561_o ? s_data : n9579_o;
  assign n9581_o = gprbit[31:24];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9582_o = n9562_o ? s_data : n9581_o;
  assign n9583_o = gprbit[39:32];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9584_o = n9563_o ? s_data : n9583_o;
  assign n9585_o = gprbit[47:40];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9586_o = n9564_o ? s_data : n9585_o;
  assign n9587_o = gprbit[55:48];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9588_o = n9565_o ? s_data : n9587_o;
  assign n9589_o = gprbit[63:56];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9590_o = n9566_o ? s_data : n9589_o;
  assign n9591_o = gprbit[71:64];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9592_o = n9567_o ? s_data : n9591_o;
  assign n9593_o = gprbit[79:72];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9594_o = n9568_o ? s_data : n9593_o;
  assign n9595_o = gprbit[87:80];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9596_o = n9569_o ? s_data : n9595_o;
  assign n9597_o = gprbit[95:88];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9598_o = n9570_o ? s_data : n9597_o;
  assign n9599_o = gprbit[103:96];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9600_o = n9571_o ? s_data : n9599_o;
  assign n9601_o = gprbit[111:104];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9602_o = n9572_o ? s_data : n9601_o;
  assign n9603_o = gprbit[119:112];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9604_o = n9573_o ? s_data : n9603_o;
  assign n9605_o = gprbit[127:120];
  /* control_mem_rtl.vhd:1059:15  */
  assign n9606_o = n9574_o ? s_data : n9605_o;
  assign n9607_o = {n9606_o, n9604_o, n9602_o, n9600_o, n9598_o, n9596_o, n9594_o, n9592_o, n9590_o, n9588_o, n9586_o, n9584_o, n9582_o, n9580_o, n9578_o, n9576_o};
  /* control_mem_rtl.vhd:1089:21  */
  assign n9608_o = n8618_o[2];
  /* control_mem_rtl.vhd:1089:21  */
  assign n9609_o = ~n9608_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9610_o = n8618_o[1];
  /* control_mem_rtl.vhd:1089:21  */
  assign n9611_o = ~n9610_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9612_o = n9609_o & n9611_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9613_o = n9609_o & n9610_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9614_o = n9608_o & n9611_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9615_o = n9608_o & n9610_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9616_o = n8618_o[0];
  /* control_mem_rtl.vhd:1089:21  */
  assign n9617_o = ~n9616_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9618_o = n9612_o & n9617_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9619_o = n9612_o & n9616_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9620_o = n9613_o & n9617_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9621_o = n9613_o & n9616_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9622_o = n9614_o & n9617_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9623_o = n9614_o & n9616_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9624_o = n9615_o & n9617_o;
  /* control_mem_rtl.vhd:1089:21  */
  assign n9625_o = n9615_o & n9616_o;
  assign n9626_o = p0[0];
  /* control_mem_rtl.vhd:1089:21  */
  assign n9627_o = n9618_o ? s_bdata : n9626_o;
  assign n9628_o = p0[1];
  /* control_mem_rtl.vhd:1089:21  */
  assign n9629_o = n9619_o ? s_bdata : n9628_o;
  assign n9630_o = p0[2];
  /* control_mem_rtl.vhd:1089:21  */
  assign n9631_o = n9620_o ? s_bdata : n9630_o;
  assign n9632_o = p0[3];
  /* control_mem_rtl.vhd:1089:21  */
  assign n9633_o = n9621_o ? s_bdata : n9632_o;
  assign n9634_o = p0[4];
  /* control_mem_rtl.vhd:1089:21  */
  assign n9635_o = n9622_o ? s_bdata : n9634_o;
  assign n9636_o = p0[5];
  /* control_mem_rtl.vhd:1089:21  */
  assign n9637_o = n9623_o ? s_bdata : n9636_o;
  assign n9638_o = p0[6];
  /* control_mem_rtl.vhd:1089:21  */
  assign n9639_o = n9624_o ? s_bdata : n9638_o;
  assign n9640_o = p0[7];
  /* control_mem_rtl.vhd:1089:21  */
  assign n9641_o = n9625_o ? s_bdata : n9640_o;
  assign n9642_o = {n9641_o, n9639_o, n9637_o, n9635_o, n9633_o, n9631_o, n9629_o, n9627_o};
  /* control_mem_rtl.vhd:1091:21  */
  assign n9643_o = n8624_o[2];
  /* control_mem_rtl.vhd:1091:21  */
  assign n9644_o = ~n9643_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9645_o = n8624_o[1];
  /* control_mem_rtl.vhd:1091:21  */
  assign n9646_o = ~n9645_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9647_o = n9644_o & n9646_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9648_o = n9644_o & n9645_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9649_o = n9643_o & n9646_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9650_o = n9643_o & n9645_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9651_o = n8624_o[0];
  /* control_mem_rtl.vhd:1091:21  */
  assign n9652_o = ~n9651_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9653_o = n9647_o & n9652_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9654_o = n9647_o & n9651_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9655_o = n9648_o & n9652_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9656_o = n9648_o & n9651_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9657_o = n9649_o & n9652_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9658_o = n9649_o & n9651_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9659_o = n9650_o & n9652_o;
  /* control_mem_rtl.vhd:1091:21  */
  assign n9660_o = n9650_o & n9651_o;
  assign n9661_o = n8631_o[0];
  /* control_mem_rtl.vhd:1091:21  */
  assign n9662_o = n9653_o ? s_bdata : n9661_o;
  assign n9663_o = n8631_o[1];
  /* control_mem_rtl.vhd:1091:21  */
  assign n9664_o = n9654_o ? s_bdata : n9663_o;
  assign n9665_o = n8631_o[2];
  /* control_mem_rtl.vhd:1091:21  */
  assign n9666_o = n9655_o ? s_bdata : n9665_o;
  assign n9667_o = n8631_o[3];
  /* control_mem_rtl.vhd:1091:21  */
  assign n9668_o = n9656_o ? s_bdata : n9667_o;
  assign n9669_o = n8631_o[4];
  /* control_mem_rtl.vhd:1091:21  */
  assign n9670_o = n9657_o ? s_bdata : n9669_o;
  assign n9671_o = n8631_o[5];
  /* control_mem_rtl.vhd:1091:21  */
  assign n9672_o = n9658_o ? s_bdata : n9671_o;
  assign n9673_o = n8631_o[6];
  /* control_mem_rtl.vhd:1091:21  */
  assign n9674_o = n9659_o ? s_bdata : n9673_o;
  assign n9675_o = n8631_o[7];
  /* control_mem_rtl.vhd:1091:21  */
  assign n9676_o = n9660_o ? s_bdata : n9675_o;
  assign n9677_o = {n9676_o, n9674_o, n9672_o, n9670_o, n9668_o, n9666_o, n9664_o, n9662_o};
  /* control_mem_rtl.vhd:1093:21  */
  assign n9678_o = n8635_o[2];
  /* control_mem_rtl.vhd:1093:21  */
  assign n9679_o = ~n9678_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9680_o = n8635_o[1];
  /* control_mem_rtl.vhd:1093:21  */
  assign n9681_o = ~n9680_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9682_o = n9679_o & n9681_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9683_o = n9679_o & n9680_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9684_o = n9678_o & n9681_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9685_o = n9678_o & n9680_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9686_o = n8635_o[0];
  /* control_mem_rtl.vhd:1093:21  */
  assign n9687_o = ~n9686_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9688_o = n9682_o & n9687_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9689_o = n9682_o & n9686_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9690_o = n9683_o & n9687_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9691_o = n9683_o & n9686_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9692_o = n9684_o & n9687_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9693_o = n9684_o & n9686_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9694_o = n9685_o & n9687_o;
  /* control_mem_rtl.vhd:1093:21  */
  assign n9695_o = n9685_o & n9686_o;
  assign n9696_o = p1[0];
  /* control_mem_rtl.vhd:1093:21  */
  assign n9697_o = n9688_o ? s_bdata : n9696_o;
  assign n9698_o = p1[1];
  /* control_mem_rtl.vhd:1093:21  */
  assign n9699_o = n9689_o ? s_bdata : n9698_o;
  assign n9700_o = p1[2];
  /* control_mem_rtl.vhd:1093:21  */
  assign n9701_o = n9690_o ? s_bdata : n9700_o;
  assign n9702_o = p1[3];
  /* control_mem_rtl.vhd:1093:21  */
  assign n9703_o = n9691_o ? s_bdata : n9702_o;
  assign n9704_o = p1[4];
  /* control_mem_rtl.vhd:1093:21  */
  assign n9705_o = n9692_o ? s_bdata : n9704_o;
  assign n9706_o = p1[5];
  /* control_mem_rtl.vhd:1093:21  */
  assign n9707_o = n9693_o ? s_bdata : n9706_o;
  assign n9708_o = p1[6];
  /* control_mem_rtl.vhd:1093:21  */
  assign n9709_o = n9694_o ? s_bdata : n9708_o;
  assign n9710_o = p1[7];
  /* control_mem_rtl.vhd:1093:21  */
  assign n9711_o = n9695_o ? s_bdata : n9710_o;
  assign n9712_o = {n9711_o, n9709_o, n9707_o, n9705_o, n9703_o, n9701_o, n9699_o, n9697_o};
  /* control_mem_rtl.vhd:1095:21  */
  assign n9713_o = n8641_o[2];
  /* control_mem_rtl.vhd:1095:21  */
  assign n9714_o = ~n9713_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9715_o = n8641_o[1];
  /* control_mem_rtl.vhd:1095:21  */
  assign n9716_o = ~n9715_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9717_o = n9714_o & n9716_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9718_o = n9714_o & n9715_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9719_o = n9713_o & n9716_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9720_o = n9713_o & n9715_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9721_o = n8641_o[0];
  /* control_mem_rtl.vhd:1095:21  */
  assign n9722_o = ~n9721_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9723_o = n9717_o & n9722_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9724_o = n9717_o & n9721_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9725_o = n9718_o & n9722_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9726_o = n9718_o & n9721_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9727_o = n9719_o & n9722_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9728_o = n9719_o & n9721_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9729_o = n9720_o & n9722_o;
  /* control_mem_rtl.vhd:1095:21  */
  assign n9730_o = n9720_o & n9721_o;
  assign n9731_o = n8645_o[0];
  /* control_mem_rtl.vhd:1095:21  */
  assign n9732_o = n9723_o ? s_bdata : n9731_o;
  assign n9733_o = n8645_o[1];
  /* control_mem_rtl.vhd:1095:21  */
  assign n9734_o = n9724_o ? s_bdata : n9733_o;
  assign n9735_o = n8645_o[2];
  /* control_mem_rtl.vhd:1095:21  */
  assign n9736_o = n9725_o ? s_bdata : n9735_o;
  assign n9737_o = n8645_o[3];
  /* control_mem_rtl.vhd:1095:21  */
  assign n9738_o = n9726_o ? s_bdata : n9737_o;
  assign n9739_o = n8645_o[4];
  /* control_mem_rtl.vhd:1095:21  */
  assign n9740_o = n9727_o ? s_bdata : n9739_o;
  assign n9741_o = n8645_o[5];
  /* control_mem_rtl.vhd:1095:21  */
  assign n9742_o = n9728_o ? s_bdata : n9741_o;
  assign n9743_o = n8645_o[6];
  /* control_mem_rtl.vhd:1095:21  */
  assign n9744_o = n9729_o ? s_bdata : n9743_o;
  assign n9745_o = n8645_o[7];
  /* control_mem_rtl.vhd:1095:21  */
  assign n9746_o = n9730_o ? s_bdata : n9745_o;
  assign n9747_o = {n9746_o, n9744_o, n9742_o, n9740_o, n9738_o, n9736_o, n9734_o, n9732_o};
  /* control_mem_rtl.vhd:1097:21  */
  assign n9748_o = n8649_o[2];
  /* control_mem_rtl.vhd:1097:21  */
  assign n9749_o = ~n9748_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9750_o = n8649_o[1];
  /* control_mem_rtl.vhd:1097:21  */
  assign n9751_o = ~n9750_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9752_o = n9749_o & n9751_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9753_o = n9749_o & n9750_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9754_o = n9748_o & n9751_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9755_o = n9748_o & n9750_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9756_o = n8649_o[0];
  /* control_mem_rtl.vhd:1097:21  */
  assign n9757_o = ~n9756_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9758_o = n9752_o & n9757_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9759_o = n9752_o & n9756_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9760_o = n9753_o & n9757_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9761_o = n9753_o & n9756_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9762_o = n9754_o & n9757_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9763_o = n9754_o & n9756_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9764_o = n9755_o & n9757_o;
  /* control_mem_rtl.vhd:1097:21  */
  assign n9765_o = n9755_o & n9756_o;
  assign n9766_o = p2[0];
  /* control_mem_rtl.vhd:1097:21  */
  assign n9767_o = n9758_o ? s_bdata : n9766_o;
  assign n9768_o = p2[1];
  /* control_mem_rtl.vhd:1097:21  */
  assign n9769_o = n9759_o ? s_bdata : n9768_o;
  assign n9770_o = p2[2];
  /* control_mem_rtl.vhd:1097:21  */
  assign n9771_o = n9760_o ? s_bdata : n9770_o;
  assign n9772_o = p2[3];
  /* control_mem_rtl.vhd:1097:21  */
  assign n9773_o = n9761_o ? s_bdata : n9772_o;
  assign n9774_o = p2[4];
  /* control_mem_rtl.vhd:1097:21  */
  assign n9775_o = n9762_o ? s_bdata : n9774_o;
  assign n9776_o = p2[5];
  /* control_mem_rtl.vhd:1097:21  */
  assign n9777_o = n9763_o ? s_bdata : n9776_o;
  assign n9778_o = p2[6];
  /* control_mem_rtl.vhd:1097:21  */
  assign n9779_o = n9764_o ? s_bdata : n9778_o;
  assign n9780_o = p2[7];
  /* control_mem_rtl.vhd:1097:21  */
  assign n9781_o = n9765_o ? s_bdata : n9780_o;
  assign n9782_o = {n9781_o, n9779_o, n9777_o, n9775_o, n9773_o, n9771_o, n9769_o, n9767_o};
  /* control_mem_rtl.vhd:1099:21  */
  assign n9783_o = n8655_o[2];
  /* control_mem_rtl.vhd:1099:21  */
  assign n9784_o = ~n9783_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9785_o = n8655_o[1];
  /* control_mem_rtl.vhd:1099:21  */
  assign n9786_o = ~n9785_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9787_o = n9784_o & n9786_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9788_o = n9784_o & n9785_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9789_o = n9783_o & n9786_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9790_o = n9783_o & n9785_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9791_o = n8655_o[0];
  /* control_mem_rtl.vhd:1099:21  */
  assign n9792_o = ~n9791_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9793_o = n9787_o & n9792_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9794_o = n9787_o & n9791_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9795_o = n9788_o & n9792_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9796_o = n9788_o & n9791_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9797_o = n9789_o & n9792_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9798_o = n9789_o & n9791_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9799_o = n9790_o & n9792_o;
  /* control_mem_rtl.vhd:1099:21  */
  assign n9800_o = n9790_o & n9791_o;
  assign n9801_o = ie[0];
  /* control_mem_rtl.vhd:1099:21  */
  assign n9802_o = n9793_o ? s_bdata : n9801_o;
  assign n9803_o = ie[1];
  /* control_mem_rtl.vhd:1099:21  */
  assign n9804_o = n9794_o ? s_bdata : n9803_o;
  assign n9805_o = ie[2];
  /* control_mem_rtl.vhd:1099:21  */
  assign n9806_o = n9795_o ? s_bdata : n9805_o;
  assign n9807_o = ie[3];
  /* control_mem_rtl.vhd:1099:21  */
  assign n9808_o = n9796_o ? s_bdata : n9807_o;
  assign n9809_o = ie[4];
  /* control_mem_rtl.vhd:1099:21  */
  assign n9810_o = n9797_o ? s_bdata : n9809_o;
  assign n9811_o = ie[5];
  /* control_mem_rtl.vhd:1099:21  */
  assign n9812_o = n9798_o ? s_bdata : n9811_o;
  assign n9813_o = ie[6];
  /* control_mem_rtl.vhd:1099:21  */
  assign n9814_o = n9799_o ? s_bdata : n9813_o;
  assign n9815_o = ie[7];
  /* control_mem_rtl.vhd:1099:21  */
  assign n9816_o = n9800_o ? s_bdata : n9815_o;
  assign n9817_o = {n9816_o, n9814_o, n9812_o, n9810_o, n9808_o, n9806_o, n9804_o, n9802_o};
  /* control_mem_rtl.vhd:1101:21  */
  assign n9818_o = n8661_o[2];
  /* control_mem_rtl.vhd:1101:21  */
  assign n9819_o = ~n9818_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9820_o = n8661_o[1];
  /* control_mem_rtl.vhd:1101:21  */
  assign n9821_o = ~n9820_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9822_o = n9819_o & n9821_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9823_o = n9819_o & n9820_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9824_o = n9818_o & n9821_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9825_o = n9818_o & n9820_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9826_o = n8661_o[0];
  /* control_mem_rtl.vhd:1101:21  */
  assign n9827_o = ~n9826_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9828_o = n9822_o & n9827_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9829_o = n9822_o & n9826_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9830_o = n9823_o & n9827_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9831_o = n9823_o & n9826_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9832_o = n9824_o & n9827_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9833_o = n9824_o & n9826_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9834_o = n9825_o & n9827_o;
  /* control_mem_rtl.vhd:1101:21  */
  assign n9835_o = n9825_o & n9826_o;
  assign n9836_o = p3[0];
  /* control_mem_rtl.vhd:1101:21  */
  assign n9837_o = n9828_o ? s_bdata : n9836_o;
  assign n9838_o = p3[1];
  /* control_mem_rtl.vhd:1101:21  */
  assign n9839_o = n9829_o ? s_bdata : n9838_o;
  assign n9840_o = p3[2];
  /* control_mem_rtl.vhd:1101:21  */
  assign n9841_o = n9830_o ? s_bdata : n9840_o;
  assign n9842_o = p3[3];
  /* control_mem_rtl.vhd:1101:21  */
  assign n9843_o = n9831_o ? s_bdata : n9842_o;
  assign n9844_o = p3[4];
  /* control_mem_rtl.vhd:1101:21  */
  assign n9845_o = n9832_o ? s_bdata : n9844_o;
  assign n9846_o = p3[5];
  /* control_mem_rtl.vhd:1101:21  */
  assign n9847_o = n9833_o ? s_bdata : n9846_o;
  assign n9848_o = p3[6];
  /* control_mem_rtl.vhd:1101:21  */
  assign n9849_o = n9834_o ? s_bdata : n9848_o;
  assign n9850_o = p3[7];
  /* control_mem_rtl.vhd:1101:21  */
  assign n9851_o = n9835_o ? s_bdata : n9850_o;
  assign n9852_o = {n9851_o, n9849_o, n9847_o, n9845_o, n9843_o, n9841_o, n9839_o, n9837_o};
  /* control_mem_rtl.vhd:1103:21  */
  assign n9853_o = n8667_o[2];
  /* control_mem_rtl.vhd:1103:21  */
  assign n9854_o = ~n9853_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9855_o = n8667_o[1];
  /* control_mem_rtl.vhd:1103:21  */
  assign n9856_o = ~n9855_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9857_o = n9854_o & n9856_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9858_o = n9854_o & n9855_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9859_o = n9853_o & n9856_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9860_o = n9853_o & n9855_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9861_o = n8667_o[0];
  /* control_mem_rtl.vhd:1103:21  */
  assign n9862_o = ~n9861_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9863_o = n9857_o & n9862_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9864_o = n9857_o & n9861_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9865_o = n9858_o & n9862_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9866_o = n9858_o & n9861_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9867_o = n9859_o & n9862_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9868_o = n9859_o & n9861_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9869_o = n9860_o & n9862_o;
  /* control_mem_rtl.vhd:1103:21  */
  assign n9870_o = n9860_o & n9861_o;
  assign n9871_o = ip[0];
  /* control_mem_rtl.vhd:1103:21  */
  assign n9872_o = n9863_o ? s_bdata : n9871_o;
  assign n9873_o = ip[1];
  /* control_mem_rtl.vhd:1103:21  */
  assign n9874_o = n9864_o ? s_bdata : n9873_o;
  assign n9875_o = ip[2];
  /* control_mem_rtl.vhd:1103:21  */
  assign n9876_o = n9865_o ? s_bdata : n9875_o;
  assign n9877_o = ip[3];
  /* control_mem_rtl.vhd:1103:21  */
  assign n9878_o = n9866_o ? s_bdata : n9877_o;
  assign n9879_o = ip[4];
  /* control_mem_rtl.vhd:1103:21  */
  assign n9880_o = n9867_o ? s_bdata : n9879_o;
  assign n9881_o = ip[5];
  /* control_mem_rtl.vhd:1103:21  */
  assign n9882_o = n9868_o ? s_bdata : n9881_o;
  assign n9883_o = ip[6];
  /* control_mem_rtl.vhd:1103:21  */
  assign n9884_o = n9869_o ? s_bdata : n9883_o;
  assign n9885_o = ip[7];
  /* control_mem_rtl.vhd:1103:21  */
  assign n9886_o = n9870_o ? s_bdata : n9885_o;
  assign n9887_o = {n9886_o, n9884_o, n9882_o, n9880_o, n9878_o, n9876_o, n9874_o, n9872_o};
  /* control_mem_rtl.vhd:1117:21  */
  assign n9888_o = n8707_o[2];
  /* control_mem_rtl.vhd:1117:21  */
  assign n9889_o = ~n9888_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9890_o = n8707_o[1];
  /* control_mem_rtl.vhd:1117:21  */
  assign n9891_o = ~n9890_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9892_o = n9889_o & n9891_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9893_o = n9889_o & n9890_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9894_o = n9888_o & n9891_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9895_o = n9888_o & n9890_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9896_o = n8707_o[0];
  /* control_mem_rtl.vhd:1117:21  */
  assign n9897_o = ~n9896_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9898_o = n9892_o & n9897_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9899_o = n9892_o & n9896_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9900_o = n9893_o & n9897_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9901_o = n9893_o & n9896_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9902_o = n9894_o & n9897_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9903_o = n9894_o & n9896_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9904_o = n9895_o & n9897_o;
  /* control_mem_rtl.vhd:1117:21  */
  assign n9905_o = n9895_o & n9896_o;
  assign n9906_o = acc[0];
  /* control_mem_rtl.vhd:1117:21  */
  assign n9907_o = n9898_o ? s_bdata : n9906_o;
  assign n9908_o = acc[1];
  /* control_mem_rtl.vhd:1117:21  */
  assign n9909_o = n9899_o ? s_bdata : n9908_o;
  assign n9910_o = acc[2];
  /* control_mem_rtl.vhd:1117:21  */
  assign n9911_o = n9900_o ? s_bdata : n9910_o;
  assign n9912_o = acc[3];
  /* control_mem_rtl.vhd:1117:21  */
  assign n9913_o = n9901_o ? s_bdata : n9912_o;
  assign n9914_o = acc[4];
  /* control_mem_rtl.vhd:1117:21  */
  assign n9915_o = n9902_o ? s_bdata : n9914_o;
  assign n9916_o = acc[5];
  /* control_mem_rtl.vhd:1117:21  */
  assign n9917_o = n9903_o ? s_bdata : n9916_o;
  assign n9918_o = acc[6];
  /* control_mem_rtl.vhd:1117:21  */
  assign n9919_o = n9904_o ? s_bdata : n9918_o;
  assign n9920_o = acc[7];
  /* control_mem_rtl.vhd:1117:21  */
  assign n9921_o = n9905_o ? s_bdata : n9920_o;
  assign n9922_o = {n9921_o, n9919_o, n9917_o, n9915_o, n9913_o, n9911_o, n9909_o, n9907_o};
  /* control_mem_rtl.vhd:1119:21  */
  assign n9923_o = n8713_o[2];
  /* control_mem_rtl.vhd:1119:21  */
  assign n9924_o = ~n9923_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9925_o = n8713_o[1];
  /* control_mem_rtl.vhd:1119:21  */
  assign n9926_o = ~n9925_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9927_o = n9924_o & n9926_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9928_o = n9924_o & n9925_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9929_o = n9923_o & n9926_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9930_o = n9923_o & n9925_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9931_o = n8713_o[0];
  /* control_mem_rtl.vhd:1119:21  */
  assign n9932_o = ~n9931_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9933_o = n9927_o & n9932_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9934_o = n9927_o & n9931_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9935_o = n9928_o & n9932_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9936_o = n9928_o & n9931_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9937_o = n9929_o & n9932_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9938_o = n9929_o & n9931_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9939_o = n9930_o & n9932_o;
  /* control_mem_rtl.vhd:1119:21  */
  assign n9940_o = n9930_o & n9931_o;
  assign n9941_o = b[0];
  /* control_mem_rtl.vhd:1119:21  */
  assign n9942_o = n9933_o ? s_bdata : n9941_o;
  assign n9943_o = b[1];
  /* control_mem_rtl.vhd:1119:21  */
  assign n9944_o = n9934_o ? s_bdata : n9943_o;
  assign n9945_o = b[2];
  /* control_mem_rtl.vhd:1119:21  */
  assign n9946_o = n9935_o ? s_bdata : n9945_o;
  assign n9947_o = b[3];
  /* control_mem_rtl.vhd:1119:21  */
  assign n9948_o = n9936_o ? s_bdata : n9947_o;
  assign n9949_o = b[4];
  /* control_mem_rtl.vhd:1119:21  */
  assign n9950_o = n9937_o ? s_bdata : n9949_o;
  assign n9951_o = b[5];
  /* control_mem_rtl.vhd:1119:21  */
  assign n9952_o = n9938_o ? s_bdata : n9951_o;
  assign n9953_o = b[6];
  /* control_mem_rtl.vhd:1119:21  */
  assign n9954_o = n9939_o ? s_bdata : n9953_o;
  assign n9955_o = b[7];
  /* control_mem_rtl.vhd:1119:21  */
  assign n9956_o = n9940_o ? s_bdata : n9955_o;
  assign n9957_o = {n9956_o, n9954_o, n9952_o, n9950_o, n9948_o, n9946_o, n9944_o, n9942_o};
  /* control_mem_rtl.vhd:1124:23  */
  assign n9958_o = {n8751_o, n8754_o};
  /* control_mem_rtl.vhd:1123:17  */
  assign n9959_o = n9958_o[6];
  /* control_mem_rtl.vhd:1123:17  */
  assign n9960_o = ~n9959_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9961_o = n9958_o[5];
  /* control_mem_rtl.vhd:1123:17  */
  assign n9962_o = ~n9961_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9963_o = n9960_o & n9962_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9964_o = n9960_o & n9961_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9965_o = n9959_o & n9962_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9966_o = n9959_o & n9961_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9967_o = n9958_o[4];
  /* control_mem_rtl.vhd:1123:17  */
  assign n9968_o = ~n9967_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9969_o = n9963_o & n9968_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9970_o = n9963_o & n9967_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9971_o = n9964_o & n9968_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9972_o = n9964_o & n9967_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9973_o = n9965_o & n9968_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9974_o = n9965_o & n9967_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9975_o = n9966_o & n9968_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9976_o = n9966_o & n9967_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9977_o = n9958_o[3];
  /* control_mem_rtl.vhd:1123:17  */
  assign n9978_o = ~n9977_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9979_o = n9969_o & n9978_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9980_o = n9969_o & n9977_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9981_o = n9970_o & n9978_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9982_o = n9970_o & n9977_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9983_o = n9971_o & n9978_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9984_o = n9971_o & n9977_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9985_o = n9972_o & n9978_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9986_o = n9972_o & n9977_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9987_o = n9973_o & n9978_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9988_o = n9973_o & n9977_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9989_o = n9974_o & n9978_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9990_o = n9974_o & n9977_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9991_o = n9975_o & n9978_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9992_o = n9975_o & n9977_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9993_o = n9976_o & n9978_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9994_o = n9976_o & n9977_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9995_o = n9958_o[2];
  /* control_mem_rtl.vhd:1123:17  */
  assign n9996_o = ~n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9997_o = n9979_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9998_o = n9979_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n9999_o = n9980_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10000_o = n9980_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10001_o = n9981_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10002_o = n9981_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10003_o = n9982_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10004_o = n9982_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10005_o = n9983_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10006_o = n9983_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10007_o = n9984_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10008_o = n9984_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10009_o = n9985_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10010_o = n9985_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10011_o = n9986_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10012_o = n9986_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10013_o = n9987_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10014_o = n9987_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10015_o = n9988_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10016_o = n9988_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10017_o = n9989_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10018_o = n9989_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10019_o = n9990_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10020_o = n9990_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10021_o = n9991_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10022_o = n9991_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10023_o = n9992_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10024_o = n9992_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10025_o = n9993_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10026_o = n9993_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10027_o = n9994_o & n9996_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10028_o = n9994_o & n9995_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10029_o = n9958_o[1];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10030_o = ~n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10031_o = n9997_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10032_o = n9997_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10033_o = n9998_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10034_o = n9998_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10035_o = n9999_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10036_o = n9999_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10037_o = n10000_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10038_o = n10000_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10039_o = n10001_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10040_o = n10001_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10041_o = n10002_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10042_o = n10002_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10043_o = n10003_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10044_o = n10003_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10045_o = n10004_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10046_o = n10004_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10047_o = n10005_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10048_o = n10005_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10049_o = n10006_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10050_o = n10006_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10051_o = n10007_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10052_o = n10007_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10053_o = n10008_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10054_o = n10008_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10055_o = n10009_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10056_o = n10009_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10057_o = n10010_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10058_o = n10010_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10059_o = n10011_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10060_o = n10011_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10061_o = n10012_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10062_o = n10012_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10063_o = n10013_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10064_o = n10013_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10065_o = n10014_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10066_o = n10014_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10067_o = n10015_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10068_o = n10015_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10069_o = n10016_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10070_o = n10016_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10071_o = n10017_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10072_o = n10017_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10073_o = n10018_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10074_o = n10018_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10075_o = n10019_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10076_o = n10019_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10077_o = n10020_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10078_o = n10020_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10079_o = n10021_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10080_o = n10021_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10081_o = n10022_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10082_o = n10022_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10083_o = n10023_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10084_o = n10023_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10085_o = n10024_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10086_o = n10024_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10087_o = n10025_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10088_o = n10025_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10089_o = n10026_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10090_o = n10026_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10091_o = n10027_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10092_o = n10027_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10093_o = n10028_o & n10030_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10094_o = n10028_o & n10029_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10095_o = n9958_o[0];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10096_o = ~n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10097_o = n10031_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10098_o = n10031_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10099_o = n10032_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10100_o = n10032_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10101_o = n10033_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10102_o = n10033_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10103_o = n10034_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10104_o = n10034_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10105_o = n10035_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10106_o = n10035_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10107_o = n10036_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10108_o = n10036_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10109_o = n10037_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10110_o = n10037_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10111_o = n10038_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10112_o = n10038_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10113_o = n10039_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10114_o = n10039_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10115_o = n10040_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10116_o = n10040_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10117_o = n10041_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10118_o = n10041_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10119_o = n10042_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10120_o = n10042_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10121_o = n10043_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10122_o = n10043_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10123_o = n10044_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10124_o = n10044_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10125_o = n10045_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10126_o = n10045_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10127_o = n10046_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10128_o = n10046_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10129_o = n10047_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10130_o = n10047_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10131_o = n10048_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10132_o = n10048_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10133_o = n10049_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10134_o = n10049_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10135_o = n10050_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10136_o = n10050_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10137_o = n10051_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10138_o = n10051_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10139_o = n10052_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10140_o = n10052_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10141_o = n10053_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10142_o = n10053_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10143_o = n10054_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10144_o = n10054_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10145_o = n10055_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10146_o = n10055_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10147_o = n10056_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10148_o = n10056_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10149_o = n10057_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10150_o = n10057_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10151_o = n10058_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10152_o = n10058_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10153_o = n10059_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10154_o = n10059_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10155_o = n10060_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10156_o = n10060_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10157_o = n10061_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10158_o = n10061_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10159_o = n10062_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10160_o = n10062_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10161_o = n10063_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10162_o = n10063_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10163_o = n10064_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10164_o = n10064_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10165_o = n10065_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10166_o = n10065_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10167_o = n10066_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10168_o = n10066_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10169_o = n10067_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10170_o = n10067_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10171_o = n10068_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10172_o = n10068_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10173_o = n10069_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10174_o = n10069_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10175_o = n10070_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10176_o = n10070_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10177_o = n10071_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10178_o = n10071_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10179_o = n10072_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10180_o = n10072_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10181_o = n10073_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10182_o = n10073_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10183_o = n10074_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10184_o = n10074_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10185_o = n10075_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10186_o = n10075_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10187_o = n10076_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10188_o = n10076_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10189_o = n10077_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10190_o = n10077_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10191_o = n10078_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10192_o = n10078_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10193_o = n10079_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10194_o = n10079_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10195_o = n10080_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10196_o = n10080_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10197_o = n10081_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10198_o = n10081_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10199_o = n10082_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10200_o = n10082_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10201_o = n10083_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10202_o = n10083_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10203_o = n10084_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10204_o = n10084_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10205_o = n10085_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10206_o = n10085_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10207_o = n10086_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10208_o = n10086_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10209_o = n10087_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10210_o = n10087_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10211_o = n10088_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10212_o = n10088_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10213_o = n10089_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10214_o = n10089_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10215_o = n10090_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10216_o = n10090_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10217_o = n10091_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10218_o = n10091_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10219_o = n10092_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10220_o = n10092_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10221_o = n10093_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10222_o = n10093_o & n10095_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10223_o = n10094_o & n10096_o;
  /* control_mem_rtl.vhd:1123:17  */
  assign n10224_o = n10094_o & n10095_o;
  assign n10225_o = gprbit[0];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10226_o = n10097_o ? s_bdata : n10225_o;
  assign n10227_o = gprbit[1];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10228_o = n10098_o ? s_bdata : n10227_o;
  assign n10229_o = gprbit[2];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10230_o = n10099_o ? s_bdata : n10229_o;
  assign n10231_o = gprbit[3];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10232_o = n10100_o ? s_bdata : n10231_o;
  assign n10233_o = gprbit[4];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10234_o = n10101_o ? s_bdata : n10233_o;
  assign n10235_o = gprbit[5];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10236_o = n10102_o ? s_bdata : n10235_o;
  assign n10237_o = gprbit[6];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10238_o = n10103_o ? s_bdata : n10237_o;
  assign n10239_o = gprbit[7];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10240_o = n10104_o ? s_bdata : n10239_o;
  assign n10241_o = gprbit[8];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10242_o = n10105_o ? s_bdata : n10241_o;
  assign n10243_o = gprbit[9];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10244_o = n10106_o ? s_bdata : n10243_o;
  assign n10245_o = gprbit[10];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10246_o = n10107_o ? s_bdata : n10245_o;
  assign n10247_o = gprbit[11];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10248_o = n10108_o ? s_bdata : n10247_o;
  assign n10249_o = gprbit[12];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10250_o = n10109_o ? s_bdata : n10249_o;
  assign n10251_o = gprbit[13];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10252_o = n10110_o ? s_bdata : n10251_o;
  assign n10253_o = gprbit[14];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10254_o = n10111_o ? s_bdata : n10253_o;
  assign n10255_o = gprbit[15];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10256_o = n10112_o ? s_bdata : n10255_o;
  assign n10257_o = gprbit[16];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10258_o = n10113_o ? s_bdata : n10257_o;
  assign n10259_o = gprbit[17];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10260_o = n10114_o ? s_bdata : n10259_o;
  assign n10261_o = gprbit[18];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10262_o = n10115_o ? s_bdata : n10261_o;
  assign n10263_o = gprbit[19];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10264_o = n10116_o ? s_bdata : n10263_o;
  assign n10265_o = gprbit[20];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10266_o = n10117_o ? s_bdata : n10265_o;
  assign n10267_o = gprbit[21];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10268_o = n10118_o ? s_bdata : n10267_o;
  assign n10269_o = gprbit[22];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10270_o = n10119_o ? s_bdata : n10269_o;
  assign n10271_o = gprbit[23];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10272_o = n10120_o ? s_bdata : n10271_o;
  assign n10273_o = gprbit[24];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10274_o = n10121_o ? s_bdata : n10273_o;
  assign n10275_o = gprbit[25];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10276_o = n10122_o ? s_bdata : n10275_o;
  assign n10277_o = gprbit[26];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10278_o = n10123_o ? s_bdata : n10277_o;
  assign n10279_o = gprbit[27];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10280_o = n10124_o ? s_bdata : n10279_o;
  assign n10281_o = gprbit[28];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10282_o = n10125_o ? s_bdata : n10281_o;
  assign n10283_o = gprbit[29];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10284_o = n10126_o ? s_bdata : n10283_o;
  assign n10285_o = gprbit[30];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10286_o = n10127_o ? s_bdata : n10285_o;
  assign n10287_o = gprbit[31];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10288_o = n10128_o ? s_bdata : n10287_o;
  assign n10289_o = gprbit[32];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10290_o = n10129_o ? s_bdata : n10289_o;
  assign n10291_o = gprbit[33];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10292_o = n10130_o ? s_bdata : n10291_o;
  assign n10293_o = gprbit[34];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10294_o = n10131_o ? s_bdata : n10293_o;
  assign n10295_o = gprbit[35];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10296_o = n10132_o ? s_bdata : n10295_o;
  assign n10297_o = gprbit[36];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10298_o = n10133_o ? s_bdata : n10297_o;
  assign n10299_o = gprbit[37];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10300_o = n10134_o ? s_bdata : n10299_o;
  assign n10301_o = gprbit[38];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10302_o = n10135_o ? s_bdata : n10301_o;
  assign n10303_o = gprbit[39];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10304_o = n10136_o ? s_bdata : n10303_o;
  assign n10305_o = gprbit[40];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10306_o = n10137_o ? s_bdata : n10305_o;
  assign n10307_o = gprbit[41];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10308_o = n10138_o ? s_bdata : n10307_o;
  assign n10309_o = gprbit[42];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10310_o = n10139_o ? s_bdata : n10309_o;
  assign n10311_o = gprbit[43];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10312_o = n10140_o ? s_bdata : n10311_o;
  assign n10313_o = gprbit[44];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10314_o = n10141_o ? s_bdata : n10313_o;
  assign n10315_o = gprbit[45];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10316_o = n10142_o ? s_bdata : n10315_o;
  assign n10317_o = gprbit[46];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10318_o = n10143_o ? s_bdata : n10317_o;
  assign n10319_o = gprbit[47];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10320_o = n10144_o ? s_bdata : n10319_o;
  assign n10321_o = gprbit[48];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10322_o = n10145_o ? s_bdata : n10321_o;
  assign n10323_o = gprbit[49];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10324_o = n10146_o ? s_bdata : n10323_o;
  assign n10325_o = gprbit[50];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10326_o = n10147_o ? s_bdata : n10325_o;
  assign n10327_o = gprbit[51];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10328_o = n10148_o ? s_bdata : n10327_o;
  assign n10329_o = gprbit[52];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10330_o = n10149_o ? s_bdata : n10329_o;
  assign n10331_o = gprbit[53];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10332_o = n10150_o ? s_bdata : n10331_o;
  assign n10333_o = gprbit[54];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10334_o = n10151_o ? s_bdata : n10333_o;
  assign n10335_o = gprbit[55];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10336_o = n10152_o ? s_bdata : n10335_o;
  assign n10337_o = gprbit[56];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10338_o = n10153_o ? s_bdata : n10337_o;
  assign n10339_o = gprbit[57];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10340_o = n10154_o ? s_bdata : n10339_o;
  assign n10341_o = gprbit[58];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10342_o = n10155_o ? s_bdata : n10341_o;
  assign n10343_o = gprbit[59];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10344_o = n10156_o ? s_bdata : n10343_o;
  assign n10345_o = gprbit[60];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10346_o = n10157_o ? s_bdata : n10345_o;
  assign n10347_o = gprbit[61];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10348_o = n10158_o ? s_bdata : n10347_o;
  assign n10349_o = gprbit[62];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10350_o = n10159_o ? s_bdata : n10349_o;
  assign n10351_o = gprbit[63];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10352_o = n10160_o ? s_bdata : n10351_o;
  assign n10353_o = gprbit[64];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10354_o = n10161_o ? s_bdata : n10353_o;
  assign n10355_o = gprbit[65];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10356_o = n10162_o ? s_bdata : n10355_o;
  assign n10357_o = gprbit[66];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10358_o = n10163_o ? s_bdata : n10357_o;
  assign n10359_o = gprbit[67];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10360_o = n10164_o ? s_bdata : n10359_o;
  assign n10361_o = gprbit[68];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10362_o = n10165_o ? s_bdata : n10361_o;
  assign n10363_o = gprbit[69];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10364_o = n10166_o ? s_bdata : n10363_o;
  assign n10365_o = gprbit[70];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10366_o = n10167_o ? s_bdata : n10365_o;
  assign n10367_o = gprbit[71];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10368_o = n10168_o ? s_bdata : n10367_o;
  assign n10369_o = gprbit[72];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10370_o = n10169_o ? s_bdata : n10369_o;
  assign n10371_o = gprbit[73];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10372_o = n10170_o ? s_bdata : n10371_o;
  assign n10373_o = gprbit[74];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10374_o = n10171_o ? s_bdata : n10373_o;
  assign n10375_o = gprbit[75];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10376_o = n10172_o ? s_bdata : n10375_o;
  assign n10377_o = gprbit[76];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10378_o = n10173_o ? s_bdata : n10377_o;
  assign n10379_o = gprbit[77];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10380_o = n10174_o ? s_bdata : n10379_o;
  assign n10381_o = gprbit[78];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10382_o = n10175_o ? s_bdata : n10381_o;
  assign n10383_o = gprbit[79];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10384_o = n10176_o ? s_bdata : n10383_o;
  assign n10385_o = gprbit[80];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10386_o = n10177_o ? s_bdata : n10385_o;
  assign n10387_o = gprbit[81];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10388_o = n10178_o ? s_bdata : n10387_o;
  assign n10389_o = gprbit[82];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10390_o = n10179_o ? s_bdata : n10389_o;
  assign n10391_o = gprbit[83];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10392_o = n10180_o ? s_bdata : n10391_o;
  assign n10393_o = gprbit[84];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10394_o = n10181_o ? s_bdata : n10393_o;
  assign n10395_o = gprbit[85];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10396_o = n10182_o ? s_bdata : n10395_o;
  assign n10397_o = gprbit[86];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10398_o = n10183_o ? s_bdata : n10397_o;
  assign n10399_o = gprbit[87];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10400_o = n10184_o ? s_bdata : n10399_o;
  assign n10401_o = gprbit[88];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10402_o = n10185_o ? s_bdata : n10401_o;
  assign n10403_o = gprbit[89];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10404_o = n10186_o ? s_bdata : n10403_o;
  assign n10405_o = gprbit[90];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10406_o = n10187_o ? s_bdata : n10405_o;
  assign n10407_o = gprbit[91];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10408_o = n10188_o ? s_bdata : n10407_o;
  assign n10409_o = gprbit[92];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10410_o = n10189_o ? s_bdata : n10409_o;
  assign n10411_o = gprbit[93];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10412_o = n10190_o ? s_bdata : n10411_o;
  assign n10413_o = gprbit[94];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10414_o = n10191_o ? s_bdata : n10413_o;
  assign n10415_o = gprbit[95];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10416_o = n10192_o ? s_bdata : n10415_o;
  assign n10417_o = gprbit[96];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10418_o = n10193_o ? s_bdata : n10417_o;
  assign n10419_o = gprbit[97];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10420_o = n10194_o ? s_bdata : n10419_o;
  assign n10421_o = gprbit[98];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10422_o = n10195_o ? s_bdata : n10421_o;
  assign n10423_o = gprbit[99];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10424_o = n10196_o ? s_bdata : n10423_o;
  assign n10425_o = gprbit[100];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10426_o = n10197_o ? s_bdata : n10425_o;
  assign n10427_o = gprbit[101];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10428_o = n10198_o ? s_bdata : n10427_o;
  assign n10429_o = gprbit[102];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10430_o = n10199_o ? s_bdata : n10429_o;
  assign n10431_o = gprbit[103];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10432_o = n10200_o ? s_bdata : n10431_o;
  assign n10433_o = gprbit[104];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10434_o = n10201_o ? s_bdata : n10433_o;
  assign n10435_o = gprbit[105];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10436_o = n10202_o ? s_bdata : n10435_o;
  assign n10437_o = gprbit[106];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10438_o = n10203_o ? s_bdata : n10437_o;
  assign n10439_o = gprbit[107];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10440_o = n10204_o ? s_bdata : n10439_o;
  assign n10441_o = gprbit[108];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10442_o = n10205_o ? s_bdata : n10441_o;
  assign n10443_o = gprbit[109];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10444_o = n10206_o ? s_bdata : n10443_o;
  assign n10445_o = gprbit[110];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10446_o = n10207_o ? s_bdata : n10445_o;
  assign n10447_o = gprbit[111];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10448_o = n10208_o ? s_bdata : n10447_o;
  assign n10449_o = gprbit[112];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10450_o = n10209_o ? s_bdata : n10449_o;
  assign n10451_o = gprbit[113];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10452_o = n10210_o ? s_bdata : n10451_o;
  assign n10453_o = gprbit[114];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10454_o = n10211_o ? s_bdata : n10453_o;
  assign n10455_o = gprbit[115];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10456_o = n10212_o ? s_bdata : n10455_o;
  assign n10457_o = gprbit[116];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10458_o = n10213_o ? s_bdata : n10457_o;
  assign n10459_o = gprbit[117];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10460_o = n10214_o ? s_bdata : n10459_o;
  assign n10461_o = gprbit[118];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10462_o = n10215_o ? s_bdata : n10461_o;
  assign n10463_o = gprbit[119];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10464_o = n10216_o ? s_bdata : n10463_o;
  assign n10465_o = gprbit[120];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10466_o = n10217_o ? s_bdata : n10465_o;
  assign n10467_o = gprbit[121];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10468_o = n10218_o ? s_bdata : n10467_o;
  assign n10469_o = gprbit[122];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10470_o = n10219_o ? s_bdata : n10469_o;
  assign n10471_o = gprbit[123];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10472_o = n10220_o ? s_bdata : n10471_o;
  assign n10473_o = gprbit[124];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10474_o = n10221_o ? s_bdata : n10473_o;
  assign n10475_o = gprbit[125];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10476_o = n10222_o ? s_bdata : n10475_o;
  assign n10477_o = gprbit[126];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10478_o = n10223_o ? s_bdata : n10477_o;
  assign n10479_o = gprbit[127];
  /* control_mem_rtl.vhd:1123:17  */
  assign n10480_o = n10224_o ? s_bdata : n10479_o;
  assign n10481_o = {n10480_o, n10478_o, n10476_o, n10474_o, n10472_o, n10470_o, n10468_o, n10466_o, n10464_o, n10462_o, n10460_o, n10458_o, n10456_o, n10454_o, n10452_o, n10450_o, n10448_o, n10446_o, n10444_o, n10442_o, n10440_o, n10438_o, n10436_o, n10434_o, n10432_o, n10430_o, n10428_o, n10426_o, n10424_o, n10422_o, n10420_o, n10418_o, n10416_o, n10414_o, n10412_o, n10410_o, n10408_o, n10406_o, n10404_o, n10402_o, n10400_o, n10398_o, n10396_o, n10394_o, n10392_o, n10390_o, n10388_o, n10386_o, n10384_o, n10382_o, n10380_o, n10378_o, n10376_o, n10374_o, n10372_o, n10370_o, n10368_o, n10366_o, n10364_o, n10362_o, n10360_o, n10358_o, n10356_o, n10354_o, n10352_o, n10350_o, n10348_o, n10346_o, n10344_o, n10342_o, n10340_o, n10338_o, n10336_o, n10334_o, n10332_o, n10330_o, n10328_o, n10326_o, n10324_o, n10322_o, n10320_o, n10318_o, n10316_o, n10314_o, n10312_o, n10310_o, n10308_o, n10306_o, n10304_o, n10302_o, n10300_o, n10298_o, n10296_o, n10294_o, n10292_o, n10290_o, n10288_o, n10286_o, n10284_o, n10282_o, n10280_o, n10278_o, n10276_o, n10274_o, n10272_o, n10270_o, n10268_o, n10266_o, n10264_o, n10262_o, n10260_o, n10258_o, n10256_o, n10254_o, n10252_o, n10250_o, n10248_o, n10246_o, n10244_o, n10242_o, n10240_o, n10238_o, n10236_o, n10234_o, n10232_o, n10230_o, n10228_o, n10226_o};
endmodule

module control_fsm
  (input  [2:0] state_i,
   input  [7:0] help_i,
   input  bit_data_i,
   input  [7:0] aludata_i,
   input  [7:0] command_i,
   input  inthigh_i,
   input  intlow_i,
   input  intpre_i,
   input  intpre2_i,
   input  intblock_i,
   input  ti_i,
   input  ri_i,
   input  ie0_i,
   input  ie1_i,
   input  tf0_i,
   input  tf1_i,
   input  [7:0] acc,
   input  [7:0] psw,
   input  [7:0] ie,
   input  [7:0] ip,
   output [5:0] alu_cmd_o,
   output [3:0] pc_inc_en_o,
   output [2:0] nextstate_o,
   output [3:0] adr_mux_o,
   output [1:0] adrx_mux_o,
   output wrx_mux_o,
   output [3:0] data_mux_o,
   output [3:0] bdata_mux_o,
   output [2:0] regs_wr_en_o,
   output [3:0] help_en_o,
   output [1:0] help16_en_o,
   output helpb_en_o,
   output inthigh_en_o,
   output intlow_en_o,
   output intpre2_en_o,
   output inthigh_d_o,
   output intlow_d_o,
   output intpre2_d_o,
   output ext0isr_d_o,
   output ext1isr_d_o,
   output ext0isrh_d_o,
   output ext1isrh_d_o,
   output ext0isr_en_o,
   output ext1isr_en_o,
   output ext0isrh_en_o,
   output ext1isrh_en_o);
  wire n2628_o;
  wire n2632_o;
  wire n2633_o;
  wire n2634_o;
  wire n2635_o;
  wire n2636_o;
  wire n2637_o;
  wire n2638_o;
  wire n2639_o;
  wire n2640_o;
  wire n2641_o;
  wire [2:0] state;
  wire [2:0] s_nextstate;
  wire [6:0] s_instr_category;
  wire [7:0] s_help;
  wire s_bit_data;
  wire s_intpre;
  wire s_intpre2;
  wire s_inthigh;
  wire s_intlow;
  wire s_tf1;
  wire s_tf0;
  wire s_ie1;
  wire s_ie0;
  wire s_ri;
  wire s_ti;
  wire [7:0] s_command;
  wire [3:0] s_pc_inc_en;
  wire [2:0] s_regs_wr_en;
  wire [3:0] s_data_mux;
  wire [3:0] s_bdata_mux;
  wire [3:0] s_adr_mux;
  wire [1:0] s_adrx_mux;
  wire s_wrx_mux;
  wire [3:0] s_help_en;
  wire [1:0] s_help16_en;
  wire s_helpb_en;
  wire s_intpre2_d;
  wire s_intpre2_en;
  wire s_intlow_d;
  wire s_intlow_en;
  wire s_inthigh_d;
  wire s_inthigh_en;
  wire s_ext0isr_d;
  wire s_ext1isr_d;
  wire s_ext0isrh_d;
  wire s_ext1isrh_d;
  wire s_ext0isr_en;
  wire s_ext1isr_en;
  wire s_ext0isrh_en;
  wire s_ext1isrh_en;
  wire [4:0] n2643_o;
  wire n2645_o;
  wire [6:0] n2646_o;
  wire [4:0] n2648_o;
  wire n2650_o;
  wire [6:0] n2651_o;
  wire n2654_o;
  wire [6:0] n2655_o;
  wire [6:0] n2657_o;
  wire n2659_o;
  wire [6:0] n2660_o;
  wire n2663_o;
  wire [6:0] n2664_o;
  wire [4:0] n2666_o;
  wire n2668_o;
  wire [6:0] n2669_o;
  wire n2672_o;
  wire [6:0] n2673_o;
  wire [6:0] n2675_o;
  wire n2677_o;
  wire [6:0] n2678_o;
  wire n2681_o;
  wire [6:0] n2682_o;
  wire [4:0] n2684_o;
  wire n2686_o;
  wire [6:0] n2687_o;
  wire [4:0] n2689_o;
  wire n2691_o;
  wire [6:0] n2692_o;
  wire n2695_o;
  wire [6:0] n2696_o;
  wire [6:0] n2698_o;
  wire n2700_o;
  wire [6:0] n2701_o;
  wire n2704_o;
  wire [6:0] n2705_o;
  wire n2708_o;
  wire [6:0] n2709_o;
  wire n2712_o;
  wire [6:0] n2713_o;
  wire n2716_o;
  wire [6:0] n2717_o;
  wire n2720_o;
  wire [6:0] n2721_o;
  wire n2724_o;
  wire [6:0] n2725_o;
  wire n2728_o;
  wire [6:0] n2729_o;
  wire [4:0] n2731_o;
  wire n2733_o;
  wire [6:0] n2734_o;
  wire [6:0] n2736_o;
  wire n2738_o;
  wire [6:0] n2739_o;
  wire n2742_o;
  wire [6:0] n2743_o;
  wire n2746_o;
  wire [6:0] n2747_o;
  wire n2750_o;
  wire [6:0] n2751_o;
  wire n2754_o;
  wire [6:0] n2755_o;
  wire n2758_o;
  wire [6:0] n2759_o;
  wire n2762_o;
  wire [6:0] n2763_o;
  wire n2766_o;
  wire [6:0] n2767_o;
  wire n2770_o;
  wire [6:0] n2771_o;
  wire [4:0] n2773_o;
  wire n2775_o;
  wire [6:0] n2776_o;
  wire n2779_o;
  wire [6:0] n2780_o;
  wire [6:0] n2782_o;
  wire n2784_o;
  wire [6:0] n2785_o;
  wire n2788_o;
  wire [6:0] n2789_o;
  wire [4:0] n2791_o;
  wire n2793_o;
  wire [6:0] n2794_o;
  wire n2797_o;
  wire [6:0] n2798_o;
  wire n2801_o;
  wire [6:0] n2802_o;
  wire [4:0] n2804_o;
  wire n2806_o;
  wire [6:0] n2807_o;
  wire n2810_o;
  wire [6:0] n2811_o;
  wire [6:0] n2813_o;
  wire n2815_o;
  wire [6:0] n2816_o;
  wire n2819_o;
  wire [6:0] n2820_o;
  wire n2823_o;
  wire [6:0] n2824_o;
  wire n2827_o;
  wire [6:0] n2828_o;
  wire n2831_o;
  wire [6:0] n2832_o;
  wire n2835_o;
  wire [6:0] n2836_o;
  wire n2839_o;
  wire [6:0] n2840_o;
  wire n2843_o;
  wire [6:0] n2844_o;
  wire n2847_o;
  wire [6:0] n2848_o;
  wire n2851_o;
  wire [6:0] n2852_o;
  wire n2855_o;
  wire [6:0] n2856_o;
  wire n2859_o;
  wire [6:0] n2860_o;
  wire [4:0] n2862_o;
  wire n2864_o;
  wire [6:0] n2865_o;
  wire n2868_o;
  wire [6:0] n2869_o;
  wire [6:0] n2871_o;
  wire n2873_o;
  wire [6:0] n2874_o;
  wire n2877_o;
  wire [6:0] n2878_o;
  wire [4:0] n2880_o;
  wire n2882_o;
  wire [6:0] n2883_o;
  wire [4:0] n2885_o;
  wire n2887_o;
  wire [6:0] n2888_o;
  wire [4:0] n2890_o;
  wire n2892_o;
  wire [6:0] n2893_o;
  wire n2896_o;
  wire [6:0] n2897_o;
  wire [4:0] n2899_o;
  wire n2901_o;
  wire [6:0] n2902_o;
  wire n2905_o;
  wire [6:0] n2906_o;
  wire [6:0] n2908_o;
  wire n2910_o;
  wire [6:0] n2911_o;
  wire n2914_o;
  wire [6:0] n2915_o;
  wire [6:0] n2917_o;
  wire n2919_o;
  wire [6:0] n2920_o;
  wire [6:0] n2922_o;
  wire n2924_o;
  wire [6:0] n2925_o;
  wire [6:0] n2927_o;
  wire n2929_o;
  wire [6:0] n2930_o;
  wire n2933_o;
  wire [6:0] n2934_o;
  wire n2937_o;
  wire [6:0] n2938_o;
  wire [6:0] n2940_o;
  wire n2942_o;
  wire [6:0] n2943_o;
  wire n2946_o;
  wire [6:0] n2947_o;
  wire [6:0] n2949_o;
  wire n2951_o;
  wire [6:0] n2952_o;
  wire n2955_o;
  wire [6:0] n2956_o;
  wire n2959_o;
  wire [6:0] n2960_o;
  wire n2963_o;
  wire [6:0] n2964_o;
  wire n2967_o;
  wire [6:0] n2968_o;
  wire n2971_o;
  wire [6:0] n2972_o;
  wire n2975_o;
  wire [6:0] n2976_o;
  wire [4:0] n2978_o;
  wire n2980_o;
  wire [6:0] n2981_o;
  wire n2984_o;
  wire [6:0] n2985_o;
  wire [6:0] n2987_o;
  wire n2989_o;
  wire [6:0] n2990_o;
  wire n2993_o;
  wire [6:0] n2994_o;
  wire n2997_o;
  wire [6:0] n2998_o;
  wire n3001_o;
  wire [6:0] n3002_o;
  wire n3005_o;
  wire [6:0] n3006_o;
  wire n3009_o;
  wire [6:0] n3010_o;
  wire n3013_o;
  wire [6:0] n3014_o;
  wire n3017_o;
  wire [6:0] n3018_o;
  wire n3021_o;
  wire [6:0] n3022_o;
  wire n3025_o;
  wire [6:0] n3026_o;
  wire n3029_o;
  wire [6:0] n3030_o;
  wire n3033_o;
  wire [6:0] n3034_o;
  wire n3037_o;
  wire [6:0] n3038_o;
  wire n3041_o;
  wire [6:0] n3042_o;
  wire n3045_o;
  wire [6:0] n3046_o;
  wire n3049_o;
  wire [6:0] n3050_o;
  wire n3053_o;
  wire [6:0] n3054_o;
  wire [4:0] n3056_o;
  wire n3058_o;
  wire [6:0] n3059_o;
  wire n3062_o;
  wire [6:0] n3063_o;
  wire [6:0] n3065_o;
  wire n3067_o;
  wire [6:0] n3068_o;
  wire n3071_o;
  wire [6:0] n3072_o;
  wire n3075_o;
  wire [6:0] n3076_o;
  wire [4:0] n3078_o;
  wire n3080_o;
  wire [6:0] n3081_o;
  wire n3084_o;
  wire [6:0] n3085_o;
  wire [6:0] n3087_o;
  wire n3089_o;
  wire [6:0] n3090_o;
  wire [6:0] n3092_o;
  wire n3094_o;
  wire [6:0] n3095_o;
  wire [4:0] n3097_o;
  wire n3099_o;
  wire [6:0] n3100_o;
  wire n3103_o;
  wire [6:0] n3104_o;
  wire [6:0] n3106_o;
  wire n3108_o;
  wire [6:0] n3109_o;
  wire n3112_o;
  wire [6:0] n3113_o;
  wire n3116_o;
  wire [6:0] n3117_o;
  wire n3120_o;
  wire [6:0] n3121_o;
  wire n3125_o;
  wire n3126_o;
  wire n3128_o;
  wire n3129_o;
  wire n3131_o;
  wire n3132_o;
  wire n3133_o;
  wire n3134_o;
  wire n3136_o;
  wire n3138_o;
  wire n3139_o;
  wire n3140_o;
  wire n3141_o;
  wire n3142_o;
  wire n3143_o;
  wire n3144_o;
  wire n3145_o;
  wire n3146_o;
  wire n3147_o;
  wire n3148_o;
  wire n3149_o;
  wire n3150_o;
  wire n3151_o;
  wire n3152_o;
  wire n3153_o;
  wire n3154_o;
  wire n3155_o;
  wire [3:0] n3158_o;
  wire n3161_o;
  wire n3164_o;
  wire [2:0] n3167_o;
  wire [3:0] n3170_o;
  wire [3:0] n3172_o;
  wire n3174_o;
  wire n3176_o;
  wire [2:0] n3178_o;
  wire [3:0] n3180_o;
  wire [3:0] n3182_o;
  wire n3184_o;
  wire n3186_o;
  wire n3189_o;
  wire n3192_o;
  wire [2:0] n3194_o;
  wire [3:0] n3196_o;
  wire [3:0] n3198_o;
  wire n3200_o;
  wire n3202_o;
  wire n3204_o;
  wire n3206_o;
  wire [2:0] n3208_o;
  wire [3:0] n3210_o;
  wire [3:0] n3212_o;
  wire n3214_o;
  wire n3216_o;
  wire n3219_o;
  wire n3221_o;
  wire n3224_o;
  wire n3226_o;
  wire [2:0] n3228_o;
  wire [3:0] n3230_o;
  wire [3:0] n3232_o;
  wire n3234_o;
  wire n3236_o;
  wire n3239_o;
  wire n3242_o;
  wire n3244_o;
  wire n3246_o;
  wire n3248_o;
  wire n3250_o;
  wire [2:0] n3252_o;
  wire [3:0] n3254_o;
  wire [3:0] n3256_o;
  wire n3258_o;
  wire n3260_o;
  wire n3262_o;
  wire n3264_o;
  wire n3266_o;
  wire n3268_o;
  wire n3270_o;
  wire n3272_o;
  wire [2:0] n3274_o;
  wire [3:0] n3276_o;
  wire [3:0] n3278_o;
  wire n3280_o;
  wire n3282_o;
  wire n3284_o;
  wire n3286_o;
  wire n3288_o;
  wire n3290_o;
  wire n3293_o;
  wire n3295_o;
  wire n3297_o;
  wire n3300_o;
  wire [2:0] n3302_o;
  wire [3:0] n3304_o;
  wire [3:0] n3306_o;
  wire n3308_o;
  wire n3310_o;
  wire n3312_o;
  wire n3314_o;
  wire n3316_o;
  wire n3318_o;
  wire n3320_o;
  wire n3322_o;
  wire n3324_o;
  wire n3326_o;
  wire [2:0] n3328_o;
  wire [3:0] n3330_o;
  wire [3:0] n3332_o;
  wire n3334_o;
  wire n3336_o;
  wire n3338_o;
  wire n3340_o;
  wire n3342_o;
  wire n3344_o;
  wire n3347_o;
  wire n3349_o;
  wire n3351_o;
  wire n3353_o;
  wire n3356_o;
  wire n3358_o;
  wire n3360_o;
  wire n3362_o;
  wire [3:0] n3365_o;
  wire [2:0] n3368_o;
  wire [3:0] n3371_o;
  wire [3:0] n3374_o;
  wire n3377_o;
  wire [2:0] n3380_o;
  wire [3:0] n3382_o;
  wire [2:0] n3384_o;
  wire [3:0] n3386_o;
  wire [3:0] n3388_o;
  wire n3390_o;
  wire [2:0] n3392_o;
  wire [3:0] n3394_o;
  wire [2:0] n3395_o;
  wire [3:0] n3397_o;
  wire [3:0] n3398_o;
  wire [3:0] n3400_o;
  wire n3402_o;
  wire n3404_o;
  wire n3406_o;
  wire n3408_o;
  wire n3410_o;
  wire n3412_o;
  wire n3414_o;
  wire n3416_o;
  wire n3418_o;
  wire n3420_o;
  wire n3422_o;
  wire n3424_o;
  wire n3426_o;
  wire [2:0] n3428_o;
  wire [3:0] n3430_o;
  wire [2:0] n3432_o;
  wire [3:0] n3434_o;
  wire [3:0] n3436_o;
  wire [3:0] n3438_o;
  wire n3441_o;
  wire n3443_o;
  wire n3445_o;
  wire n3447_o;
  wire n3449_o;
  wire n3451_o;
  wire n3453_o;
  wire n3455_o;
  wire n3457_o;
  wire n3459_o;
  wire n3461_o;
  wire n3463_o;
  wire n3465_o;
  wire n3467_o;
  wire n3469_o;
  wire n3471_o;
  wire [3:0] n3474_o;
  wire [2:0] n3477_o;
  wire [3:0] n3480_o;
  wire [3:0] n3483_o;
  wire [2:0] n3486_o;
  wire [3:0] n3488_o;
  wire [2:0] n3490_o;
  wire [3:0] n3492_o;
  wire [3:0] n3494_o;
  wire [1:0] n3497_o;
  wire n3499_o;
  wire n3501_o;
  wire n3503_o;
  wire [5:0] n3506_o;
  wire [3:0] n3509_o;
  wire [2:0] n3512_o;
  wire [3:0] n3515_o;
  wire [5:0] n3517_o;
  wire [2:0] n3520_o;
  wire [3:0] n3522_o;
  wire [2:0] n3524_o;
  wire [3:0] n3526_o;
  wire [3:0] n3529_o;
  wire n3531_o;
  wire n3533_o;
  wire n3535_o;
  wire n3537_o;
  wire [5:0] n3540_o;
  wire [3:0] n3543_o;
  wire [2:0] n3546_o;
  wire [3:0] n3549_o;
  wire [5:0] n3551_o;
  wire [2:0] n3554_o;
  wire [3:0] n3556_o;
  wire [2:0] n3558_o;
  wire [3:0] n3560_o;
  wire [3:0] n3563_o;
  wire [5:0] n3565_o;
  wire [2:0] n3567_o;
  wire [3:0] n3569_o;
  wire [2:0] n3571_o;
  wire [3:0] n3573_o;
  wire [3:0] n3575_o;
  wire n3577_o;
  wire n3579_o;
  wire n3581_o;
  wire [5:0] n3584_o;
  wire [3:0] n3587_o;
  wire [2:0] n3590_o;
  wire [3:0] n3593_o;
  wire [5:0] n3595_o;
  wire [2:0] n3598_o;
  wire [3:0] n3600_o;
  wire [2:0] n3602_o;
  wire [3:0] n3604_o;
  wire [3:0] n3607_o;
  wire n3609_o;
  wire n3611_o;
  wire n3613_o;
  wire [5:0] n3616_o;
  wire [3:0] n3619_o;
  wire [2:0] n3622_o;
  wire [3:0] n3625_o;
  wire [5:0] n3627_o;
  wire [2:0] n3630_o;
  wire [3:0] n3632_o;
  wire [2:0] n3634_o;
  wire [3:0] n3636_o;
  wire n3638_o;
  wire n3640_o;
  wire n3642_o;
  wire [5:0] n3645_o;
  wire [3:0] n3648_o;
  wire [2:0] n3651_o;
  wire [3:0] n3654_o;
  wire [5:0] n3656_o;
  wire [2:0] n3659_o;
  wire [3:0] n3661_o;
  wire [2:0] n3663_o;
  wire [3:0] n3665_o;
  wire [3:0] n3668_o;
  wire n3670_o;
  wire n3672_o;
  wire n3674_o;
  wire n3676_o;
  wire [5:0] n3679_o;
  wire [3:0] n3682_o;
  wire [2:0] n3685_o;
  wire [3:0] n3688_o;
  wire [5:0] n3690_o;
  wire [2:0] n3693_o;
  wire [3:0] n3695_o;
  wire [2:0] n3697_o;
  wire [3:0] n3699_o;
  wire [3:0] n3702_o;
  wire [5:0] n3704_o;
  wire [2:0] n3706_o;
  wire [3:0] n3708_o;
  wire [2:0] n3710_o;
  wire [3:0] n3712_o;
  wire [3:0] n3714_o;
  wire n3716_o;
  wire n3718_o;
  wire n3720_o;
  wire [5:0] n3723_o;
  wire [3:0] n3726_o;
  wire [2:0] n3729_o;
  wire [3:0] n3732_o;
  wire [5:0] n3734_o;
  wire [2:0] n3737_o;
  wire [3:0] n3739_o;
  wire [2:0] n3741_o;
  wire [3:0] n3743_o;
  wire [3:0] n3746_o;
  wire n3748_o;
  wire n3750_o;
  wire n3752_o;
  wire [5:0] n3755_o;
  wire [3:0] n3758_o;
  wire [2:0] n3761_o;
  wire [3:0] n3764_o;
  wire [5:0] n3766_o;
  wire [2:0] n3769_o;
  wire [3:0] n3771_o;
  wire [2:0] n3773_o;
  wire [3:0] n3775_o;
  wire n3777_o;
  wire n3779_o;
  wire n3781_o;
  wire [3:0] n3784_o;
  wire [2:0] n3787_o;
  wire [3:0] n3789_o;
  wire [1:0] n3792_o;
  wire n3794_o;
  wire n3796_o;
  wire n3798_o;
  wire [5:0] n3801_o;
  wire [3:0] n3804_o;
  wire [2:0] n3807_o;
  wire [3:0] n3810_o;
  wire [5:0] n3812_o;
  wire [2:0] n3815_o;
  wire [3:0] n3817_o;
  wire [2:0] n3819_o;
  wire [3:0] n3821_o;
  wire [3:0] n3824_o;
  wire n3826_o;
  wire n3828_o;
  wire n3830_o;
  wire n3832_o;
  wire [5:0] n3835_o;
  wire [3:0] n3838_o;
  wire [2:0] n3841_o;
  wire [3:0] n3844_o;
  wire [5:0] n3846_o;
  wire [2:0] n3849_o;
  wire [3:0] n3851_o;
  wire [2:0] n3853_o;
  wire [3:0] n3855_o;
  wire [3:0] n3858_o;
  wire [5:0] n3860_o;
  wire [2:0] n3862_o;
  wire [3:0] n3864_o;
  wire [2:0] n3866_o;
  wire [3:0] n3868_o;
  wire [3:0] n3870_o;
  wire n3872_o;
  wire n3874_o;
  wire n3876_o;
  wire [5:0] n3879_o;
  wire [3:0] n3882_o;
  wire [2:0] n3885_o;
  wire [3:0] n3888_o;
  wire [5:0] n3890_o;
  wire [2:0] n3893_o;
  wire [3:0] n3895_o;
  wire [2:0] n3897_o;
  wire [3:0] n3899_o;
  wire [3:0] n3902_o;
  wire n3904_o;
  wire n3906_o;
  wire n3908_o;
  wire [5:0] n3911_o;
  wire [3:0] n3914_o;
  wire [2:0] n3917_o;
  wire [3:0] n3920_o;
  wire [5:0] n3922_o;
  wire [2:0] n3925_o;
  wire [3:0] n3927_o;
  wire [2:0] n3929_o;
  wire [3:0] n3931_o;
  wire n3933_o;
  wire n3935_o;
  wire n3937_o;
  wire n3939_o;
  wire [5:0] n3942_o;
  wire [3:0] n3945_o;
  wire [2:0] n3948_o;
  wire [3:0] n3951_o;
  wire [3:0] n3954_o;
  wire [5:0] n3956_o;
  wire [2:0] n3959_o;
  wire [3:0] n3961_o;
  wire [2:0] n3963_o;
  wire [3:0] n3965_o;
  wire [3:0] n3967_o;
  wire [5:0] n3969_o;
  wire [2:0] n3971_o;
  wire [3:0] n3973_o;
  wire [2:0] n3975_o;
  wire [3:0] n3977_o;
  wire [3:0] n3979_o;
  wire n3981_o;
  wire n3983_o;
  wire n3985_o;
  wire n3987_o;
  wire [5:0] n3990_o;
  wire [3:0] n3993_o;
  wire [2:0] n3996_o;
  wire [3:0] n3999_o;
  wire [3:0] n4002_o;
  wire [5:0] n4004_o;
  wire [2:0] n4007_o;
  wire [3:0] n4009_o;
  wire [2:0] n4011_o;
  wire [3:0] n4013_o;
  wire [3:0] n4015_o;
  wire [3:0] n4018_o;
  wire [5:0] n4020_o;
  wire [2:0] n4022_o;
  wire [3:0] n4024_o;
  wire [2:0] n4026_o;
  wire [3:0] n4028_o;
  wire [3:0] n4030_o;
  wire [3:0] n4032_o;
  wire n4034_o;
  wire n4036_o;
  wire n4038_o;
  wire n4040_o;
  wire [3:0] n4043_o;
  wire [2:0] n4046_o;
  wire [3:0] n4049_o;
  wire [2:0] n4052_o;
  wire [3:0] n4054_o;
  wire [2:0] n4056_o;
  wire [3:0] n4058_o;
  wire [3:0] n4061_o;
  wire [2:0] n4063_o;
  wire [3:0] n4065_o;
  wire [2:0] n4067_o;
  wire [3:0] n4069_o;
  wire [3:0] n4071_o;
  wire n4073_o;
  wire n4075_o;
  wire n4077_o;
  wire n4079_o;
  wire [3:0] n4082_o;
  wire [2:0] n4085_o;
  wire [3:0] n4088_o;
  wire [2:0] n4091_o;
  wire [3:0] n4093_o;
  wire [2:0] n4095_o;
  wire [3:0] n4097_o;
  wire [3:0] n4100_o;
  wire [2:0] n4102_o;
  wire [3:0] n4104_o;
  wire [2:0] n4106_o;
  wire [3:0] n4108_o;
  wire [3:0] n4110_o;
  wire n4112_o;
  wire n4114_o;
  wire n4116_o;
  wire n4118_o;
  wire [8:0] n4119_o;
  wire n4121_o;
  wire [3:0] n4124_o;
  wire [3:0] n4127_o;
  wire [5:0] n4130_o;
  wire [3:0] n4132_o;
  wire [2:0] n4135_o;
  wire [3:0] n4137_o;
  wire [3:0] n4140_o;
  wire [5:0] n4142_o;
  wire [2:0] n4145_o;
  wire [3:0] n4147_o;
  wire [2:0] n4149_o;
  wire [3:0] n4151_o;
  wire [3:0] n4153_o;
  wire [5:0] n4155_o;
  wire [2:0] n4157_o;
  wire [3:0] n4159_o;
  wire [2:0] n4161_o;
  wire [3:0] n4163_o;
  wire [3:0] n4165_o;
  wire n4167_o;
  wire n4169_o;
  wire n4171_o;
  wire n4173_o;
  wire [8:0] n4174_o;
  wire n4176_o;
  wire [3:0] n4179_o;
  wire [3:0] n4182_o;
  wire [3:0] n4184_o;
  wire [2:0] n4187_o;
  wire [3:0] n4189_o;
  wire [3:0] n4192_o;
  wire [5:0] n4195_o;
  wire [2:0] n4198_o;
  wire [3:0] n4200_o;
  wire [2:0] n4202_o;
  wire [3:0] n4204_o;
  wire [3:0] n4206_o;
  wire [3:0] n4209_o;
  wire n4212_o;
  wire [5:0] n4214_o;
  wire [2:0] n4216_o;
  wire [3:0] n4218_o;
  wire [2:0] n4220_o;
  wire [3:0] n4222_o;
  wire [3:0] n4224_o;
  wire [3:0] n4226_o;
  wire n4228_o;
  wire n4230_o;
  wire n4232_o;
  wire n4234_o;
  wire n4236_o;
  wire [8:0] n4237_o;
  wire n4239_o;
  wire [3:0] n4242_o;
  wire [3:0] n4245_o;
  wire [3:0] n4247_o;
  wire [2:0] n4250_o;
  wire [3:0] n4252_o;
  wire [3:0] n4255_o;
  wire [5:0] n4258_o;
  wire [2:0] n4261_o;
  wire [3:0] n4263_o;
  wire [2:0] n4265_o;
  wire [3:0] n4267_o;
  wire [3:0] n4269_o;
  wire [3:0] n4272_o;
  wire n4275_o;
  wire [5:0] n4277_o;
  wire [2:0] n4279_o;
  wire [3:0] n4281_o;
  wire [2:0] n4283_o;
  wire [3:0] n4285_o;
  wire [3:0] n4287_o;
  wire [3:0] n4289_o;
  wire n4291_o;
  wire n4293_o;
  wire n4295_o;
  wire n4297_o;
  wire n4299_o;
  wire [8:0] n4300_o;
  wire n4302_o;
  wire [3:0] n4305_o;
  wire [3:0] n4308_o;
  wire [3:0] n4310_o;
  wire [2:0] n4313_o;
  wire [3:0] n4315_o;
  wire [3:0] n4318_o;
  wire [5:0] n4321_o;
  wire [2:0] n4324_o;
  wire [3:0] n4326_o;
  wire [2:0] n4328_o;
  wire [3:0] n4330_o;
  wire [3:0] n4332_o;
  wire [3:0] n4335_o;
  wire n4338_o;
  wire [5:0] n4340_o;
  wire [2:0] n4342_o;
  wire [3:0] n4344_o;
  wire [2:0] n4346_o;
  wire [3:0] n4348_o;
  wire [3:0] n4350_o;
  wire [3:0] n4352_o;
  wire n4354_o;
  wire n4356_o;
  wire n4358_o;
  wire n4360_o;
  wire n4362_o;
  wire n4364_o;
  wire [3:0] n4367_o;
  wire [2:0] n4370_o;
  wire [3:0] n4373_o;
  wire [2:0] n4376_o;
  wire [3:0] n4378_o;
  wire [2:0] n4380_o;
  wire [3:0] n4382_o;
  wire n4384_o;
  wire n4386_o;
  wire n4388_o;
  wire n4390_o;
  wire n4392_o;
  wire n4394_o;
  wire [3:0] n4397_o;
  wire [2:0] n4400_o;
  wire [3:0] n4403_o;
  wire [3:0] n4406_o;
  wire [2:0] n4409_o;
  wire [3:0] n4411_o;
  wire [2:0] n4413_o;
  wire [3:0] n4415_o;
  wire [3:0] n4417_o;
  wire [2:0] n4419_o;
  wire [3:0] n4421_o;
  wire [2:0] n4423_o;
  wire [3:0] n4425_o;
  wire [3:0] n4427_o;
  wire n4429_o;
  wire n4431_o;
  wire n4433_o;
  wire n4435_o;
  wire n4437_o;
  wire [5:0] n4440_o;
  wire [3:0] n4443_o;
  wire [2:0] n4446_o;
  wire [3:0] n4449_o;
  wire [3:0] n4452_o;
  wire [5:0] n4454_o;
  wire [2:0] n4457_o;
  wire [3:0] n4459_o;
  wire [2:0] n4461_o;
  wire [3:0] n4463_o;
  wire [3:0] n4465_o;
  wire n4467_o;
  wire n4469_o;
  wire n4471_o;
  wire n4473_o;
  wire [5:0] n4476_o;
  wire [3:0] n4479_o;
  wire [2:0] n4482_o;
  wire [3:0] n4485_o;
  wire [3:0] n4488_o;
  wire [5:0] n4490_o;
  wire [2:0] n4493_o;
  wire [3:0] n4495_o;
  wire [2:0] n4497_o;
  wire [3:0] n4499_o;
  wire [3:0] n4501_o;
  wire [5:0] n4503_o;
  wire [2:0] n4505_o;
  wire [3:0] n4507_o;
  wire [2:0] n4509_o;
  wire [3:0] n4511_o;
  wire [3:0] n4513_o;
  wire n4515_o;
  wire n4517_o;
  wire n4519_o;
  wire [5:0] n4522_o;
  wire [3:0] n4525_o;
  wire [2:0] n4528_o;
  wire [3:0] n4531_o;
  wire [3:0] n4534_o;
  wire [5:0] n4536_o;
  wire [2:0] n4539_o;
  wire [3:0] n4541_o;
  wire [2:0] n4543_o;
  wire [3:0] n4545_o;
  wire [3:0] n4547_o;
  wire n4549_o;
  wire n4551_o;
  wire n4553_o;
  wire n4555_o;
  wire [5:0] n4558_o;
  wire [3:0] n4561_o;
  wire [2:0] n4564_o;
  wire [3:0] n4567_o;
  wire [3:0] n4570_o;
  wire [5:0] n4572_o;
  wire [2:0] n4575_o;
  wire [3:0] n4577_o;
  wire [2:0] n4579_o;
  wire [3:0] n4581_o;
  wire [3:0] n4583_o;
  wire [5:0] n4585_o;
  wire [2:0] n4587_o;
  wire [3:0] n4589_o;
  wire [2:0] n4591_o;
  wire [3:0] n4593_o;
  wire [3:0] n4595_o;
  wire n4597_o;
  wire n4599_o;
  wire n4601_o;
  wire [8:0] n4602_o;
  wire n4604_o;
  wire [3:0] n4607_o;
  wire [5:0] n4610_o;
  wire [3:0] n4612_o;
  wire [2:0] n4615_o;
  wire [3:0] n4618_o;
  wire [3:0] n4621_o;
  wire [5:0] n4623_o;
  wire [2:0] n4626_o;
  wire [3:0] n4628_o;
  wire [2:0] n4630_o;
  wire [3:0] n4632_o;
  wire [3:0] n4634_o;
  wire [3:0] n4637_o;
  wire n4639_o;
  wire n4641_o;
  wire n4643_o;
  wire n4645_o;
  wire [8:0] n4646_o;
  wire n4648_o;
  wire [3:0] n4651_o;
  wire [5:0] n4654_o;
  wire [3:0] n4656_o;
  wire [2:0] n4659_o;
  wire [3:0] n4662_o;
  wire [3:0] n4665_o;
  wire [5:0] n4667_o;
  wire [2:0] n4670_o;
  wire [3:0] n4672_o;
  wire [2:0] n4674_o;
  wire [3:0] n4676_o;
  wire [3:0] n4678_o;
  wire [3:0] n4681_o;
  wire [5:0] n4683_o;
  wire [2:0] n4685_o;
  wire [3:0] n4687_o;
  wire [2:0] n4689_o;
  wire [3:0] n4691_o;
  wire [3:0] n4693_o;
  wire [3:0] n4695_o;
  wire n4697_o;
  wire n4699_o;
  wire n4701_o;
  wire n4703_o;
  wire [5:0] n4706_o;
  wire [3:0] n4709_o;
  wire [2:0] n4712_o;
  wire [3:0] n4715_o;
  wire [3:0] n4718_o;
  wire [5:0] n4720_o;
  wire [2:0] n4723_o;
  wire [3:0] n4725_o;
  wire [2:0] n4727_o;
  wire [3:0] n4729_o;
  wire [3:0] n4731_o;
  wire n4733_o;
  wire n4735_o;
  wire n4737_o;
  wire n4739_o;
  wire [5:0] n4742_o;
  wire [3:0] n4745_o;
  wire [2:0] n4748_o;
  wire [3:0] n4751_o;
  wire [3:0] n4754_o;
  wire [5:0] n4756_o;
  wire [2:0] n4759_o;
  wire [3:0] n4761_o;
  wire [2:0] n4763_o;
  wire [3:0] n4765_o;
  wire [3:0] n4767_o;
  wire [5:0] n4769_o;
  wire [2:0] n4771_o;
  wire [3:0] n4773_o;
  wire [2:0] n4775_o;
  wire [3:0] n4777_o;
  wire [3:0] n4779_o;
  wire n4781_o;
  wire n4783_o;
  wire n4785_o;
  wire [5:0] n4788_o;
  wire [3:0] n4791_o;
  wire [2:0] n4794_o;
  wire [3:0] n4797_o;
  wire [3:0] n4800_o;
  wire [5:0] n4802_o;
  wire [2:0] n4805_o;
  wire [3:0] n4807_o;
  wire [2:0] n4809_o;
  wire [3:0] n4811_o;
  wire [3:0] n4813_o;
  wire n4815_o;
  wire n4817_o;
  wire n4819_o;
  wire n4821_o;
  wire n4823_o;
  wire n4825_o;
  wire [5:0] n4828_o;
  wire [2:0] n4831_o;
  wire [3:0] n4834_o;
  wire [3:0] n4837_o;
  wire [5:0] n4839_o;
  wire [3:0] n4842_o;
  wire [2:0] n4844_o;
  wire [3:0] n4846_o;
  wire [3:0] n4848_o;
  wire [5:0] n4850_o;
  wire [2:0] n4853_o;
  wire [3:0] n4855_o;
  wire [2:0] n4857_o;
  wire [3:0] n4859_o;
  wire [3:0] n4861_o;
  wire [5:0] n4863_o;
  wire [2:0] n4865_o;
  wire [3:0] n4867_o;
  wire [2:0] n4869_o;
  wire [3:0] n4871_o;
  wire [3:0] n4873_o;
  wire [3:0] n4876_o;
  wire [5:0] n4878_o;
  wire [2:0] n4880_o;
  wire [3:0] n4882_o;
  wire [2:0] n4884_o;
  wire [3:0] n4886_o;
  wire [3:0] n4888_o;
  wire [3:0] n4890_o;
  wire n4892_o;
  wire n4894_o;
  wire n4896_o;
  wire n4898_o;
  wire [3:0] n4901_o;
  wire [3:0] n4903_o;
  wire [2:0] n4906_o;
  wire [3:0] n4908_o;
  wire [3:0] n4911_o;
  wire [2:0] n4913_o;
  wire [3:0] n4915_o;
  wire [3:0] n4917_o;
  wire n4919_o;
  wire n4921_o;
  wire n4923_o;
  wire n4925_o;
  wire [3:0] n4928_o;
  wire [3:0] n4930_o;
  wire [2:0] n4933_o;
  wire [3:0] n4936_o;
  wire [2:0] n4939_o;
  wire [3:0] n4941_o;
  wire [2:0] n4943_o;
  wire [3:0] n4945_o;
  wire [3:0] n4948_o;
  wire [2:0] n4950_o;
  wire [3:0] n4952_o;
  wire [2:0] n4954_o;
  wire [3:0] n4956_o;
  wire [3:0] n4958_o;
  wire n4960_o;
  wire n4962_o;
  wire n4964_o;
  wire [3:0] n4967_o;
  wire [3:0] n4969_o;
  wire [2:0] n4972_o;
  wire [3:0] n4974_o;
  wire n4976_o;
  wire n4978_o;
  wire n4980_o;
  wire n4982_o;
  wire n4984_o;
  wire n4985_o;
  wire [3:0] n4988_o;
  wire [3:0] n4990_o;
  wire [2:0] n4993_o;
  wire [3:0] n4995_o;
  wire [3:0] n4998_o;
  wire [2:0] n5000_o;
  wire [3:0] n5002_o;
  wire [3:0] n5004_o;
  wire n5006_o;
  wire n5008_o;
  wire n5010_o;
  wire n5011_o;
  wire [3:0] n5014_o;
  wire [3:0] n5016_o;
  wire [2:0] n5019_o;
  wire [3:0] n5021_o;
  wire n5023_o;
  wire n5025_o;
  wire n5027_o;
  wire n5029_o;
  wire [3:0] n5032_o;
  wire [3:0] n5034_o;
  wire [2:0] n5037_o;
  wire [3:0] n5039_o;
  wire n5041_o;
  wire n5043_o;
  wire n5045_o;
  wire n5047_o;
  wire [3:0] n5050_o;
  wire [3:0] n5052_o;
  wire [2:0] n5055_o;
  wire [3:0] n5057_o;
  wire n5059_o;
  wire n5061_o;
  wire n5063_o;
  wire n5065_o;
  wire [3:0] n5068_o;
  wire [2:0] n5071_o;
  wire [3:0] n5074_o;
  wire [3:0] n5077_o;
  wire [2:0] n5080_o;
  wire [3:0] n5082_o;
  wire [2:0] n5084_o;
  wire [3:0] n5086_o;
  wire [3:0] n5088_o;
  wire [3:0] n5091_o;
  wire [2:0] n5093_o;
  wire [3:0] n5095_o;
  wire [2:0] n5097_o;
  wire [3:0] n5099_o;
  wire [3:0] n5101_o;
  wire [3:0] n5103_o;
  wire [1:0] n5106_o;
  wire n5108_o;
  wire n5110_o;
  wire n5112_o;
  wire n5114_o;
  wire [3:0] n5117_o;
  wire [2:0] n5120_o;
  wire [3:0] n5122_o;
  wire [3:0] n5125_o;
  wire [2:0] n5127_o;
  wire [3:0] n5129_o;
  wire [3:0] n5131_o;
  wire n5133_o;
  wire n5135_o;
  wire n5137_o;
  wire [3:0] n5140_o;
  wire [2:0] n5143_o;
  wire [3:0] n5146_o;
  wire [2:0] n5149_o;
  wire [3:0] n5151_o;
  wire [2:0] n5153_o;
  wire [3:0] n5155_o;
  wire [3:0] n5158_o;
  wire n5160_o;
  wire n5162_o;
  wire n5164_o;
  wire n5166_o;
  wire [3:0] n5169_o;
  wire [2:0] n5172_o;
  wire [3:0] n5175_o;
  wire [2:0] n5178_o;
  wire [3:0] n5180_o;
  wire [2:0] n5182_o;
  wire [3:0] n5184_o;
  wire [3:0] n5187_o;
  wire [2:0] n5189_o;
  wire [3:0] n5191_o;
  wire [2:0] n5193_o;
  wire [3:0] n5195_o;
  wire [3:0] n5197_o;
  wire n5199_o;
  wire n5201_o;
  wire n5203_o;
  wire [3:0] n5206_o;
  wire [2:0] n5209_o;
  wire [3:0] n5212_o;
  wire [2:0] n5215_o;
  wire [3:0] n5217_o;
  wire [2:0] n5219_o;
  wire [3:0] n5221_o;
  wire [3:0] n5224_o;
  wire n5226_o;
  wire n5228_o;
  wire n5230_o;
  wire [3:0] n5233_o;
  wire [2:0] n5236_o;
  wire [3:0] n5239_o;
  wire [2:0] n5242_o;
  wire [3:0] n5244_o;
  wire [2:0] n5246_o;
  wire [3:0] n5248_o;
  wire n5250_o;
  wire n5252_o;
  wire n5254_o;
  wire n5256_o;
  wire n5258_o;
  wire [3:0] n5261_o;
  wire [2:0] n5264_o;
  wire [3:0] n5267_o;
  wire [3:0] n5270_o;
  wire [2:0] n5273_o;
  wire [3:0] n5275_o;
  wire [2:0] n5277_o;
  wire [3:0] n5279_o;
  wire [3:0] n5281_o;
  wire [2:0] n5283_o;
  wire [3:0] n5285_o;
  wire [2:0] n5287_o;
  wire [3:0] n5289_o;
  wire [3:0] n5291_o;
  wire [3:0] n5294_o;
  wire n5296_o;
  wire n5298_o;
  wire n5300_o;
  wire [3:0] n5303_o;
  wire [2:0] n5306_o;
  wire [3:0] n5309_o;
  wire [3:0] n5312_o;
  wire [2:0] n5315_o;
  wire [3:0] n5317_o;
  wire [2:0] n5319_o;
  wire [3:0] n5321_o;
  wire [3:0] n5323_o;
  wire [3:0] n5326_o;
  wire n5328_o;
  wire n5330_o;
  wire n5332_o;
  wire [3:0] n5335_o;
  wire [2:0] n5338_o;
  wire [3:0] n5341_o;
  wire [3:0] n5344_o;
  wire [2:0] n5347_o;
  wire [3:0] n5349_o;
  wire [2:0] n5351_o;
  wire [3:0] n5353_o;
  wire [3:0] n5355_o;
  wire n5357_o;
  wire n5359_o;
  wire n5361_o;
  wire [3:0] n5364_o;
  wire [2:0] n5367_o;
  wire [3:0] n5370_o;
  wire [3:0] n5373_o;
  wire [2:0] n5376_o;
  wire [3:0] n5378_o;
  wire [2:0] n5380_o;
  wire [3:0] n5382_o;
  wire [3:0] n5384_o;
  wire n5386_o;
  wire n5388_o;
  wire n5390_o;
  wire n5392_o;
  wire [3:0] n5395_o;
  wire [2:0] n5398_o;
  wire [3:0] n5401_o;
  wire [3:0] n5404_o;
  wire [2:0] n5407_o;
  wire [3:0] n5409_o;
  wire [2:0] n5411_o;
  wire [3:0] n5413_o;
  wire [3:0] n5415_o;
  wire [2:0] n5417_o;
  wire [3:0] n5419_o;
  wire [2:0] n5421_o;
  wire [3:0] n5423_o;
  wire [3:0] n5425_o;
  wire n5427_o;
  wire n5429_o;
  wire n5431_o;
  wire [3:0] n5434_o;
  wire [2:0] n5437_o;
  wire [3:0] n5440_o;
  wire [3:0] n5443_o;
  wire [2:0] n5446_o;
  wire [3:0] n5448_o;
  wire [2:0] n5450_o;
  wire [3:0] n5452_o;
  wire [3:0] n5454_o;
  wire n5456_o;
  wire n5458_o;
  wire n5460_o;
  wire n5462_o;
  wire [3:0] n5465_o;
  wire [2:0] n5468_o;
  wire [3:0] n5471_o;
  wire [3:0] n5474_o;
  wire [2:0] n5477_o;
  wire [3:0] n5479_o;
  wire [2:0] n5481_o;
  wire [3:0] n5483_o;
  wire [3:0] n5485_o;
  wire [3:0] n5488_o;
  wire [2:0] n5490_o;
  wire [3:0] n5492_o;
  wire [2:0] n5494_o;
  wire [3:0] n5496_o;
  wire [3:0] n5498_o;
  wire [3:0] n5500_o;
  wire n5502_o;
  wire n5504_o;
  wire n5506_o;
  wire n5508_o;
  wire n5510_o;
  wire [3:0] n5513_o;
  wire [2:0] n5516_o;
  wire [3:0] n5519_o;
  wire [3:0] n5522_o;
  wire [2:0] n5525_o;
  wire [3:0] n5527_o;
  wire [2:0] n5529_o;
  wire [3:0] n5531_o;
  wire [3:0] n5533_o;
  wire [2:0] n5535_o;
  wire [3:0] n5537_o;
  wire [2:0] n5539_o;
  wire [3:0] n5541_o;
  wire [3:0] n5543_o;
  wire n5545_o;
  wire n5547_o;
  wire n5549_o;
  wire [3:0] n5552_o;
  wire [2:0] n5555_o;
  wire [3:0] n5558_o;
  wire [3:0] n5561_o;
  wire [2:0] n5564_o;
  wire [3:0] n5566_o;
  wire [2:0] n5568_o;
  wire [3:0] n5570_o;
  wire [3:0] n5572_o;
  wire n5574_o;
  wire n5576_o;
  wire n5578_o;
  wire [3:0] n5581_o;
  wire [2:0] n5584_o;
  wire [3:0] n5587_o;
  wire [2:0] n5590_o;
  wire [3:0] n5592_o;
  wire [2:0] n5594_o;
  wire [3:0] n5596_o;
  wire [1:0] n5599_o;
  wire n5601_o;
  wire n5603_o;
  wire n5605_o;
  wire [3:0] n5608_o;
  wire [2:0] n5611_o;
  wire [3:0] n5614_o;
  wire [2:0] n5617_o;
  wire [3:0] n5619_o;
  wire [2:0] n5621_o;
  wire [3:0] n5623_o;
  wire [1:0] n5626_o;
  wire n5628_o;
  wire n5630_o;
  wire n5632_o;
  wire [3:0] n5635_o;
  wire [2:0] n5638_o;
  wire [3:0] n5641_o;
  wire [2:0] n5644_o;
  wire [3:0] n5646_o;
  wire [2:0] n5648_o;
  wire [3:0] n5650_o;
  wire [1:0] n5653_o;
  wire n5655_o;
  wire n5657_o;
  wire n5659_o;
  wire [3:0] n5662_o;
  wire [2:0] n5665_o;
  wire [3:0] n5668_o;
  wire [2:0] n5671_o;
  wire [3:0] n5673_o;
  wire [2:0] n5675_o;
  wire [3:0] n5677_o;
  wire [1:0] n5680_o;
  wire n5682_o;
  wire n5684_o;
  wire n5686_o;
  wire n5688_o;
  wire n5690_o;
  wire n5692_o;
  wire [3:0] n5695_o;
  wire [2:0] n5698_o;
  wire [3:0] n5701_o;
  wire [2:0] n5704_o;
  wire [3:0] n5706_o;
  wire [2:0] n5708_o;
  wire [3:0] n5710_o;
  wire [3:0] n5713_o;
  wire [2:0] n5715_o;
  wire [3:0] n5717_o;
  wire [2:0] n5719_o;
  wire [3:0] n5721_o;
  wire [3:0] n5723_o;
  wire n5725_o;
  wire n5727_o;
  wire n5729_o;
  wire [3:0] n5732_o;
  wire [2:0] n5735_o;
  wire [3:0] n5738_o;
  wire [3:0] n5741_o;
  wire [2:0] n5744_o;
  wire [3:0] n5746_o;
  wire [2:0] n5748_o;
  wire [3:0] n5750_o;
  wire [3:0] n5752_o;
  wire n5754_o;
  wire n5756_o;
  wire n5758_o;
  wire n5760_o;
  wire [3:0] n5763_o;
  wire [2:0] n5766_o;
  wire [3:0] n5769_o;
  wire [3:0] n5772_o;
  wire [2:0] n5775_o;
  wire [3:0] n5777_o;
  wire [2:0] n5779_o;
  wire [3:0] n5781_o;
  wire [3:0] n5783_o;
  wire [2:0] n5785_o;
  wire [3:0] n5787_o;
  wire [2:0] n5789_o;
  wire [3:0] n5791_o;
  wire [3:0] n5793_o;
  wire n5795_o;
  wire n5797_o;
  wire n5799_o;
  wire n5801_o;
  wire [5:0] n5804_o;
  wire [3:0] n5807_o;
  wire [2:0] n5810_o;
  wire [3:0] n5813_o;
  wire [3:0] n5816_o;
  wire [5:0] n5818_o;
  wire [2:0] n5821_o;
  wire [3:0] n5823_o;
  wire [2:0] n5825_o;
  wire [3:0] n5827_o;
  wire [3:0] n5829_o;
  wire [5:0] n5831_o;
  wire [2:0] n5833_o;
  wire [3:0] n5835_o;
  wire [2:0] n5837_o;
  wire [3:0] n5839_o;
  wire [3:0] n5841_o;
  wire n5843_o;
  wire n5845_o;
  wire n5847_o;
  wire n5849_o;
  wire [5:0] n5852_o;
  wire [3:0] n5855_o;
  wire [2:0] n5858_o;
  wire [3:0] n5861_o;
  wire [5:0] n5863_o;
  wire [2:0] n5866_o;
  wire [3:0] n5868_o;
  wire [2:0] n5870_o;
  wire [3:0] n5872_o;
  wire [3:0] n5875_o;
  wire n5877_o;
  wire n5879_o;
  wire n5881_o;
  wire n5883_o;
  wire [5:0] n5886_o;
  wire [3:0] n5889_o;
  wire [2:0] n5892_o;
  wire [3:0] n5895_o;
  wire [5:0] n5897_o;
  wire [2:0] n5900_o;
  wire [3:0] n5902_o;
  wire [2:0] n5904_o;
  wire [3:0] n5906_o;
  wire [3:0] n5909_o;
  wire [5:0] n5911_o;
  wire [2:0] n5913_o;
  wire [3:0] n5915_o;
  wire [2:0] n5917_o;
  wire [3:0] n5919_o;
  wire [3:0] n5921_o;
  wire n5923_o;
  wire n5925_o;
  wire n5927_o;
  wire [5:0] n5930_o;
  wire [3:0] n5933_o;
  wire [2:0] n5936_o;
  wire [3:0] n5939_o;
  wire [5:0] n5941_o;
  wire [2:0] n5944_o;
  wire [3:0] n5946_o;
  wire [2:0] n5948_o;
  wire [3:0] n5950_o;
  wire [3:0] n5953_o;
  wire n5955_o;
  wire n5957_o;
  wire n5959_o;
  wire [5:0] n5962_o;
  wire [3:0] n5965_o;
  wire [2:0] n5968_o;
  wire [3:0] n5971_o;
  wire [5:0] n5973_o;
  wire [2:0] n5976_o;
  wire [3:0] n5978_o;
  wire [2:0] n5980_o;
  wire [3:0] n5982_o;
  wire n5984_o;
  wire n5986_o;
  wire n5988_o;
  wire n5990_o;
  wire [5:0] n5993_o;
  wire [3:0] n5996_o;
  wire [2:0] n5999_o;
  wire [3:0] n6002_o;
  wire [3:0] n6005_o;
  wire [5:0] n6007_o;
  wire [2:0] n6010_o;
  wire [3:0] n6012_o;
  wire [2:0] n6014_o;
  wire [3:0] n6016_o;
  wire [3:0] n6018_o;
  wire [5:0] n6020_o;
  wire [2:0] n6022_o;
  wire [3:0] n6024_o;
  wire [2:0] n6026_o;
  wire [3:0] n6028_o;
  wire [3:0] n6030_o;
  wire n6032_o;
  wire n6034_o;
  wire n6036_o;
  wire n6038_o;
  wire [5:0] n6041_o;
  wire [3:0] n6044_o;
  wire [2:0] n6047_o;
  wire [3:0] n6050_o;
  wire [3:0] n6053_o;
  wire [5:0] n6055_o;
  wire [2:0] n6058_o;
  wire [3:0] n6060_o;
  wire [2:0] n6062_o;
  wire [3:0] n6064_o;
  wire [3:0] n6066_o;
  wire [3:0] n6069_o;
  wire [5:0] n6071_o;
  wire [2:0] n6073_o;
  wire [3:0] n6075_o;
  wire [2:0] n6077_o;
  wire [3:0] n6079_o;
  wire [3:0] n6081_o;
  wire [3:0] n6083_o;
  wire n6085_o;
  wire n6087_o;
  wire n6089_o;
  wire n6091_o;
  wire [3:0] n6094_o;
  wire [2:0] n6097_o;
  wire [3:0] n6100_o;
  wire [2:0] n6103_o;
  wire [3:0] n6105_o;
  wire [2:0] n6107_o;
  wire [3:0] n6109_o;
  wire [3:0] n6112_o;
  wire [2:0] n6114_o;
  wire [3:0] n6116_o;
  wire [2:0] n6118_o;
  wire [3:0] n6120_o;
  wire [3:0] n6122_o;
  wire n6124_o;
  wire n6126_o;
  wire n6128_o;
  wire n6130_o;
  wire [3:0] n6133_o;
  wire [2:0] n6136_o;
  wire [3:0] n6139_o;
  wire [2:0] n6142_o;
  wire [3:0] n6144_o;
  wire [2:0] n6146_o;
  wire [3:0] n6148_o;
  wire [3:0] n6151_o;
  wire [2:0] n6153_o;
  wire [3:0] n6155_o;
  wire [2:0] n6157_o;
  wire [3:0] n6159_o;
  wire [3:0] n6161_o;
  wire n6163_o;
  wire n6165_o;
  wire n6167_o;
  wire [3:0] n6170_o;
  wire [2:0] n6173_o;
  wire [3:0] n6176_o;
  wire [3:0] n6179_o;
  wire [2:0] n6182_o;
  wire [3:0] n6184_o;
  wire [2:0] n6186_o;
  wire [3:0] n6188_o;
  wire [3:0] n6190_o;
  wire n6192_o;
  wire n6194_o;
  wire n6196_o;
  wire n6198_o;
  wire [3:0] n6201_o;
  wire [2:0] n6204_o;
  wire [3:0] n6207_o;
  wire [3:0] n6210_o;
  wire [2:0] n6213_o;
  wire [3:0] n6215_o;
  wire [2:0] n6217_o;
  wire [3:0] n6219_o;
  wire [3:0] n6221_o;
  wire [2:0] n6223_o;
  wire [3:0] n6225_o;
  wire [2:0] n6227_o;
  wire [3:0] n6229_o;
  wire [3:0] n6231_o;
  wire n6233_o;
  wire n6235_o;
  wire n6237_o;
  wire n6239_o;
  wire [3:0] n6242_o;
  wire [2:0] n6245_o;
  wire [2:0] n6248_o;
  wire [3:0] n6250_o;
  wire [2:0] n6252_o;
  wire [3:0] n6255_o;
  wire [3:0] n6258_o;
  wire [2:0] n6260_o;
  wire [3:0] n6262_o;
  wire [2:0] n6264_o;
  wire [3:0] n6266_o;
  wire [3:0] n6268_o;
  wire n6270_o;
  wire n6272_o;
  wire n6274_o;
  wire n6276_o;
  wire n6279_o;
  wire n6282_o;
  wire n6285_o;
  wire n6287_o;
  wire n6290_o;
  wire n6292_o;
  wire n6294_o;
  wire n6297_o;
  wire n6300_o;
  wire [3:0] n6303_o;
  wire [2:0] n6306_o;
  wire n6308_o;
  wire n6310_o;
  wire n6312_o;
  wire n6314_o;
  wire n6316_o;
  wire n6318_o;
  wire [2:0] n6321_o;
  wire [3:0] n6323_o;
  wire [2:0] n6325_o;
  wire [3:0] n6328_o;
  wire [3:0] n6331_o;
  wire n6333_o;
  wire n6335_o;
  wire n6337_o;
  wire n6339_o;
  wire n6341_o;
  wire n6343_o;
  wire [2:0] n6345_o;
  wire [3:0] n6347_o;
  wire [2:0] n6349_o;
  wire [3:0] n6351_o;
  wire [3:0] n6353_o;
  wire n6355_o;
  wire n6357_o;
  wire n6359_o;
  wire n6361_o;
  wire n6363_o;
  wire n6365_o;
  wire n6367_o;
  wire n6369_o;
  wire n6371_o;
  wire n6373_o;
  wire n6375_o;
  wire n6377_o;
  wire n6379_o;
  wire n6381_o;
  wire [3:0] n6384_o;
  wire [2:0] n6387_o;
  wire [3:0] n6390_o;
  wire [3:0] n6393_o;
  wire [2:0] n6396_o;
  wire [3:0] n6398_o;
  wire [2:0] n6400_o;
  wire [3:0] n6402_o;
  wire [3:0] n6404_o;
  wire n6406_o;
  wire n6408_o;
  wire n6410_o;
  wire [3:0] n6413_o;
  wire [2:0] n6416_o;
  wire [3:0] n6418_o;
  wire n6420_o;
  wire n6422_o;
  wire n6424_o;
  wire [5:0] n6427_o;
  wire [3:0] n6430_o;
  wire [2:0] n6433_o;
  wire [3:0] n6436_o;
  wire [5:0] n6438_o;
  wire [2:0] n6441_o;
  wire [3:0] n6443_o;
  wire [2:0] n6445_o;
  wire [3:0] n6447_o;
  wire [3:0] n6450_o;
  wire n6452_o;
  wire n6454_o;
  wire n6456_o;
  wire n6458_o;
  wire [5:0] n6461_o;
  wire [3:0] n6464_o;
  wire [2:0] n6467_o;
  wire [3:0] n6470_o;
  wire [5:0] n6472_o;
  wire [2:0] n6475_o;
  wire [3:0] n6477_o;
  wire [2:0] n6479_o;
  wire [3:0] n6481_o;
  wire [3:0] n6484_o;
  wire [5:0] n6486_o;
  wire [2:0] n6488_o;
  wire [3:0] n6490_o;
  wire [2:0] n6492_o;
  wire [3:0] n6494_o;
  wire [3:0] n6496_o;
  wire n6498_o;
  wire n6500_o;
  wire n6502_o;
  wire [5:0] n6505_o;
  wire [3:0] n6508_o;
  wire [2:0] n6511_o;
  wire [3:0] n6514_o;
  wire [5:0] n6516_o;
  wire [2:0] n6519_o;
  wire [3:0] n6521_o;
  wire [2:0] n6523_o;
  wire [3:0] n6525_o;
  wire [3:0] n6528_o;
  wire n6530_o;
  wire n6532_o;
  wire n6534_o;
  wire [5:0] n6537_o;
  wire [3:0] n6540_o;
  wire [2:0] n6543_o;
  wire [3:0] n6546_o;
  wire [5:0] n6548_o;
  wire [2:0] n6551_o;
  wire [3:0] n6553_o;
  wire [2:0] n6555_o;
  wire [3:0] n6557_o;
  wire n6559_o;
  wire n6561_o;
  wire n6563_o;
  wire n6565_o;
  wire n6567_o;
  wire [3:0] n6570_o;
  wire [2:0] n6573_o;
  wire [3:0] n6576_o;
  wire [2:0] n6579_o;
  wire [3:0] n6581_o;
  wire [2:0] n6583_o;
  wire [3:0] n6585_o;
  wire [3:0] n6588_o;
  wire [3:0] n6591_o;
  wire [2:0] n6593_o;
  wire [3:0] n6595_o;
  wire [2:0] n6597_o;
  wire [3:0] n6599_o;
  wire [3:0] n6601_o;
  wire [3:0] n6603_o;
  wire n6605_o;
  wire n6607_o;
  wire n6609_o;
  wire n6611_o;
  wire n6613_o;
  wire [3:0] n6616_o;
  wire [2:0] n6619_o;
  wire [3:0] n6622_o;
  wire [2:0] n6625_o;
  wire [3:0] n6627_o;
  wire [2:0] n6629_o;
  wire [3:0] n6631_o;
  wire [3:0] n6634_o;
  wire [3:0] n6637_o;
  wire [2:0] n6639_o;
  wire [3:0] n6641_o;
  wire [2:0] n6643_o;
  wire [3:0] n6645_o;
  wire [3:0] n6647_o;
  wire [3:0] n6649_o;
  wire [2:0] n6651_o;
  wire [3:0] n6653_o;
  wire [2:0] n6655_o;
  wire [3:0] n6657_o;
  wire [3:0] n6659_o;
  wire [3:0] n6661_o;
  wire n6663_o;
  wire n6665_o;
  wire n6667_o;
  wire n6669_o;
  wire [3:0] n6672_o;
  wire [2:0] n6675_o;
  wire [3:0] n6678_o;
  wire [2:0] n6681_o;
  wire [3:0] n6683_o;
  wire [2:0] n6685_o;
  wire [3:0] n6687_o;
  wire [3:0] n6690_o;
  wire [3:0] n6693_o;
  wire [2:0] n6695_o;
  wire [3:0] n6697_o;
  wire [2:0] n6699_o;
  wire [3:0] n6701_o;
  wire [3:0] n6703_o;
  wire [3:0] n6705_o;
  wire n6707_o;
  wire n6709_o;
  wire n6711_o;
  wire n6713_o;
  wire [3:0] n6716_o;
  wire [2:0] n6719_o;
  wire [3:0] n6722_o;
  wire [3:0] n6725_o;
  wire [2:0] n6728_o;
  wire [3:0] n6730_o;
  wire [2:0] n6732_o;
  wire [3:0] n6734_o;
  wire [3:0] n6736_o;
  wire [2:0] n6738_o;
  wire [3:0] n6740_o;
  wire [2:0] n6742_o;
  wire [3:0] n6744_o;
  wire [3:0] n6746_o;
  wire [3:0] n6749_o;
  wire n6751_o;
  wire n6753_o;
  wire n6755_o;
  wire [5:0] n6758_o;
  wire [3:0] n6761_o;
  wire [2:0] n6764_o;
  wire [3:0] n6767_o;
  wire [5:0] n6769_o;
  wire [2:0] n6772_o;
  wire [3:0] n6774_o;
  wire [2:0] n6776_o;
  wire [3:0] n6778_o;
  wire [3:0] n6781_o;
  wire n6783_o;
  wire n6785_o;
  wire n6787_o;
  wire n6789_o;
  wire [5:0] n6792_o;
  wire [3:0] n6795_o;
  wire [2:0] n6798_o;
  wire [3:0] n6801_o;
  wire [5:0] n6803_o;
  wire [2:0] n6806_o;
  wire [3:0] n6808_o;
  wire [2:0] n6810_o;
  wire [3:0] n6812_o;
  wire [3:0] n6815_o;
  wire [5:0] n6817_o;
  wire [2:0] n6819_o;
  wire [3:0] n6821_o;
  wire [2:0] n6823_o;
  wire [3:0] n6825_o;
  wire [3:0] n6827_o;
  wire n6829_o;
  wire n6831_o;
  wire n6833_o;
  wire [5:0] n6836_o;
  wire [3:0] n6839_o;
  wire [2:0] n6842_o;
  wire [3:0] n6845_o;
  wire [5:0] n6847_o;
  wire [2:0] n6850_o;
  wire [3:0] n6852_o;
  wire [2:0] n6854_o;
  wire [3:0] n6856_o;
  wire [3:0] n6859_o;
  wire n6861_o;
  wire n6863_o;
  wire n6865_o;
  wire [5:0] n6868_o;
  wire [3:0] n6871_o;
  wire [2:0] n6874_o;
  wire [3:0] n6877_o;
  wire [5:0] n6879_o;
  wire [2:0] n6882_o;
  wire [3:0] n6884_o;
  wire [2:0] n6886_o;
  wire [3:0] n6888_o;
  wire n6890_o;
  wire n6892_o;
  wire n6894_o;
  wire n6896_o;
  wire [5:0] n6899_o;
  wire [3:0] n6902_o;
  wire [2:0] n6905_o;
  wire [3:0] n6908_o;
  wire [3:0] n6911_o;
  wire [5:0] n6913_o;
  wire [2:0] n6916_o;
  wire [3:0] n6918_o;
  wire [2:0] n6920_o;
  wire [3:0] n6922_o;
  wire [3:0] n6924_o;
  wire [5:0] n6926_o;
  wire [2:0] n6928_o;
  wire [3:0] n6930_o;
  wire [2:0] n6932_o;
  wire [3:0] n6934_o;
  wire [3:0] n6936_o;
  wire n6938_o;
  wire n6940_o;
  wire n6942_o;
  wire n6944_o;
  wire [5:0] n6947_o;
  wire [3:0] n6950_o;
  wire [2:0] n6953_o;
  wire [3:0] n6956_o;
  wire [3:0] n6959_o;
  wire [5:0] n6961_o;
  wire [2:0] n6964_o;
  wire [3:0] n6966_o;
  wire [2:0] n6968_o;
  wire [3:0] n6970_o;
  wire [3:0] n6972_o;
  wire [3:0] n6975_o;
  wire [5:0] n6977_o;
  wire [2:0] n6979_o;
  wire [3:0] n6981_o;
  wire [2:0] n6983_o;
  wire [3:0] n6985_o;
  wire [3:0] n6987_o;
  wire [3:0] n6989_o;
  wire n6991_o;
  wire [110:0] n6992_o;
  reg [5:0] n7002_o;
  reg [2:0] n7023_o;
  reg [3:0] n7044_o;
  reg [2:0] n7061_o;
  reg [3:0] n7075_o;
  reg [3:0] n7080_o;
  reg [3:0] n7087_o;
  reg [1:0] n7091_o;
  reg n7095_o;
  reg [3:0] n7097_o;
  reg [1:0] n7099_o;
  reg n7101_o;
  reg n7103_o;
  reg n7105_o;
  reg n7107_o;
  reg n7109_o;
  reg n7111_o;
  reg n7113_o;
  wire [5:0] n7115_o;
  wire [2:0] n7116_o;
  wire [3:0] n7117_o;
  wire [2:0] n7118_o;
  wire [3:0] n7119_o;
  wire [3:0] n7121_o;
  wire [3:0] n7122_o;
  wire [1:0] n7124_o;
  wire n7126_o;
  wire [3:0] n7127_o;
  wire [1:0] n7129_o;
  wire n7131_o;
  wire n7133_o;
  wire n7135_o;
  wire n7137_o;
  wire n7138_o;
  wire n7140_o;
  wire n7141_o;
  wire n7143_o;
  wire n7145_o;
  wire n7147_o;
  wire n7149_o;
  wire n7150_o;
  wire n7151_o;
  wire n7152_o;
  wire n7153_o;
  wire [5:0] n7155_o;
  wire [2:0] n7158_o;
  wire [3:0] n7161_o;
  wire [2:0] n7164_o;
  wire [3:0] n7167_o;
  wire [3:0] n7170_o;
  wire [3:0] n7173_o;
  wire [1:0] n7176_o;
  wire n7179_o;
  wire [3:0] n7182_o;
  wire [1:0] n7185_o;
  wire n7188_o;
  wire n7191_o;
  wire n7194_o;
  wire n7197_o;
  wire n7200_o;
  wire n7203_o;
  wire n7206_o;
  wire n7209_o;
  wire n7212_o;
  wire n7215_o;
  wire n7218_o;
  wire n7221_o;
  wire n7224_o;
  wire n7227_o;
  wire n7230_o;
  assign alu_cmd_o = n7155_o;
  assign pc_inc_en_o = s_pc_inc_en;
  assign nextstate_o = s_nextstate;
  assign adr_mux_o = s_adr_mux;
  assign adrx_mux_o = s_adrx_mux;
  assign wrx_mux_o = s_wrx_mux;
  assign data_mux_o = s_data_mux;
  assign bdata_mux_o = s_bdata_mux;
  assign regs_wr_en_o = s_regs_wr_en;
  assign help_en_o = s_help_en;
  assign help16_en_o = s_help16_en;
  assign helpb_en_o = s_helpb_en;
  assign inthigh_en_o = s_inthigh_en;
  assign intlow_en_o = s_intlow_en;
  assign intpre2_en_o = s_intpre2_en;
  assign inthigh_d_o = s_inthigh_d;
  assign intlow_d_o = s_intlow_d;
  assign intpre2_d_o = s_intpre2_d;
  assign ext0isr_d_o = s_ext0isr_d;
  assign ext1isr_d_o = s_ext1isr_d;
  assign ext0isrh_d_o = s_ext0isrh_d;
  assign ext1isrh_d_o = s_ext1isrh_d;
  assign ext0isr_en_o = s_ext0isr_en;
  assign ext1isr_en_o = s_ext1isr_en;
  assign ext0isrh_en_o = s_ext0isrh_en;
  assign ext1isrh_en_o = s_ext1isrh_en;
  assign n2628_o = psw[7];
  assign n2632_o = ie[4];
  /* mc8051_tmrctr_rtl.vhd:241:34  */
  assign n2633_o = ie[3];
  /* mc8051_tmrctr_rtl.vhd:226:3  */
  assign n2634_o = ie[2];
  assign n2635_o = ie[1];
  /* mc8051_tmrctr_rtl.vhd:202:9  */
  assign n2636_o = ie[0];
  /* mc8051_tmrctr_rtl.vhd:202:9  */
  assign n2637_o = ip[4];
  /* mc8051_tmrctr_rtl.vhd:202:9  */
  assign n2638_o = ip[3];
  assign n2639_o = ip[2];
  /* mc8051_tmrctr_rtl.vhd:193:3  */
  assign n2640_o = ip[1];
  assign n2641_o = ip[0];
  /* control_fsm_rtl.vhd:83:10  */
  assign state = state_i; // (signal)
  /* control_fsm_rtl.vhd:84:10  */
  assign s_nextstate = n7158_o; // (signal)
  /* control_fsm_rtl.vhd:85:10  */
  assign s_instr_category = n2646_o; // (signal)
  /* control_fsm_rtl.vhd:87:10  */
  assign s_help = help_i; // (signal)
  /* control_fsm_rtl.vhd:89:10  */
  assign s_bit_data = bit_data_i; // (signal)
  /* control_fsm_rtl.vhd:90:10  */
  assign s_intpre = intpre_i; // (signal)
  /* control_fsm_rtl.vhd:91:10  */
  assign s_intpre2 = intpre2_i; // (signal)
  /* control_fsm_rtl.vhd:92:10  */
  assign s_inthigh = inthigh_i; // (signal)
  /* control_fsm_rtl.vhd:93:10  */
  assign s_intlow = intlow_i; // (signal)
  /* control_fsm_rtl.vhd:95:10  */
  assign s_tf1 = tf1_i; // (signal)
  /* control_fsm_rtl.vhd:96:10  */
  assign s_tf0 = tf0_i; // (signal)
  /* control_fsm_rtl.vhd:97:10  */
  assign s_ie1 = ie1_i; // (signal)
  /* control_fsm_rtl.vhd:98:10  */
  assign s_ie0 = ie0_i; // (signal)
  /* control_fsm_rtl.vhd:100:10  */
  assign s_ri = ri_i; // (signal)
  /* control_fsm_rtl.vhd:101:10  */
  assign s_ti = ti_i; // (signal)
  /* control_fsm_rtl.vhd:103:10  */
  assign s_command = command_i; // (signal)
  /* control_fsm_rtl.vhd:105:10  */
  assign s_pc_inc_en = n7161_o; // (signal)
  /* control_fsm_rtl.vhd:106:10  */
  assign s_regs_wr_en = n7164_o; // (signal)
  /* control_fsm_rtl.vhd:107:10  */
  assign s_data_mux = n7167_o; // (signal)
  /* control_fsm_rtl.vhd:108:10  */
  assign s_bdata_mux = n7170_o; // (signal)
  /* control_fsm_rtl.vhd:109:10  */
  assign s_adr_mux = n7173_o; // (signal)
  /* control_fsm_rtl.vhd:110:10  */
  assign s_adrx_mux = n7176_o; // (signal)
  /* control_fsm_rtl.vhd:111:10  */
  assign s_wrx_mux = n7179_o; // (signal)
  /* control_fsm_rtl.vhd:112:10  */
  assign s_help_en = n7182_o; // (signal)
  /* control_fsm_rtl.vhd:113:10  */
  assign s_help16_en = n7185_o; // (signal)
  /* control_fsm_rtl.vhd:114:10  */
  assign s_helpb_en = n7188_o; // (signal)
  /* control_fsm_rtl.vhd:115:10  */
  assign s_intpre2_d = n7191_o; // (signal)
  /* control_fsm_rtl.vhd:116:10  */
  assign s_intpre2_en = n7194_o; // (signal)
  /* control_fsm_rtl.vhd:117:10  */
  assign s_intlow_d = n7197_o; // (signal)
  /* control_fsm_rtl.vhd:118:10  */
  assign s_intlow_en = n7200_o; // (signal)
  /* control_fsm_rtl.vhd:119:10  */
  assign s_inthigh_d = n7203_o; // (signal)
  /* control_fsm_rtl.vhd:120:10  */
  assign s_inthigh_en = n7206_o; // (signal)
  /* control_fsm_rtl.vhd:121:10  */
  assign s_ext0isr_d = n7209_o; // (signal)
  /* control_fsm_rtl.vhd:122:10  */
  assign s_ext1isr_d = n7212_o; // (signal)
  /* control_fsm_rtl.vhd:123:10  */
  assign s_ext0isrh_d = n7215_o; // (signal)
  /* control_fsm_rtl.vhd:124:10  */
  assign s_ext1isrh_d = n7218_o; // (signal)
  /* control_fsm_rtl.vhd:125:10  */
  assign s_ext0isr_en = n7221_o; // (signal)
  /* control_fsm_rtl.vhd:126:10  */
  assign s_ext1isr_en = n7224_o; // (signal)
  /* control_fsm_rtl.vhd:127:10  */
  assign s_ext0isrh_en = n7227_o; // (signal)
  /* control_fsm_rtl.vhd:128:10  */
  assign s_ext1isrh_en = n7230_o; // (signal)
  /* control_fsm_rtl.vhd:179:37  */
  assign n2643_o = s_command[4:0];
  /* control_fsm_rtl.vhd:179:50  */
  assign n2645_o = n2643_o == 5'b10001;
  /* control_fsm_rtl.vhd:179:23  */
  assign n2646_o = n2645_o ? 7'b0000000 : n2651_o;
  /* control_fsm_rtl.vhd:180:37  */
  assign n2648_o = s_command[7:3];
  /* control_fsm_rtl.vhd:180:50  */
  assign n2650_o = n2648_o == 5'b00101;
  /* control_fsm_rtl.vhd:179:67  */
  assign n2651_o = n2650_o ? 7'b0000001 : n2655_o;
  /* control_fsm_rtl.vhd:181:50  */
  assign n2654_o = s_command == 8'b00100101;
  /* control_fsm_rtl.vhd:180:67  */
  assign n2655_o = n2654_o ? 7'b0000010 : n2660_o;
  /* control_fsm_rtl.vhd:182:37  */
  assign n2657_o = s_command[7:1];
  /* control_fsm_rtl.vhd:182:50  */
  assign n2659_o = n2657_o == 7'b0010011;
  /* control_fsm_rtl.vhd:181:67  */
  assign n2660_o = n2659_o ? 7'b0000011 : n2664_o;
  /* control_fsm_rtl.vhd:183:50  */
  assign n2663_o = s_command == 8'b00100100;
  /* control_fsm_rtl.vhd:182:67  */
  assign n2664_o = n2663_o ? 7'b0000100 : n2669_o;
  /* control_fsm_rtl.vhd:184:37  */
  assign n2666_o = s_command[7:3];
  /* control_fsm_rtl.vhd:184:50  */
  assign n2668_o = n2666_o == 5'b00111;
  /* control_fsm_rtl.vhd:183:67  */
  assign n2669_o = n2668_o ? 7'b0000101 : n2673_o;
  /* control_fsm_rtl.vhd:185:50  */
  assign n2672_o = s_command == 8'b00110101;
  /* control_fsm_rtl.vhd:184:67  */
  assign n2673_o = n2672_o ? 7'b0000110 : n2678_o;
  /* control_fsm_rtl.vhd:186:37  */
  assign n2675_o = s_command[7:1];
  /* control_fsm_rtl.vhd:186:50  */
  assign n2677_o = n2675_o == 7'b0011011;
  /* control_fsm_rtl.vhd:185:67  */
  assign n2678_o = n2677_o ? 7'b0000111 : n2682_o;
  /* control_fsm_rtl.vhd:187:50  */
  assign n2681_o = s_command == 8'b00110100;
  /* control_fsm_rtl.vhd:186:67  */
  assign n2682_o = n2681_o ? 7'b0001000 : n2687_o;
  /* control_fsm_rtl.vhd:188:37  */
  assign n2684_o = s_command[4:0];
  /* control_fsm_rtl.vhd:188:50  */
  assign n2686_o = n2684_o == 5'b00001;
  /* control_fsm_rtl.vhd:187:67  */
  assign n2687_o = n2686_o ? 7'b0001001 : n2692_o;
  /* control_fsm_rtl.vhd:189:37  */
  assign n2689_o = s_command[7:3];
  /* control_fsm_rtl.vhd:189:50  */
  assign n2691_o = n2689_o == 5'b01011;
  /* control_fsm_rtl.vhd:188:67  */
  assign n2692_o = n2691_o ? 7'b0001010 : n2696_o;
  /* control_fsm_rtl.vhd:190:50  */
  assign n2695_o = s_command == 8'b01010101;
  /* control_fsm_rtl.vhd:189:67  */
  assign n2696_o = n2695_o ? 7'b0001011 : n2701_o;
  /* control_fsm_rtl.vhd:191:37  */
  assign n2698_o = s_command[7:1];
  /* control_fsm_rtl.vhd:191:50  */
  assign n2700_o = n2698_o == 7'b0101011;
  /* control_fsm_rtl.vhd:190:67  */
  assign n2701_o = n2700_o ? 7'b0001100 : n2705_o;
  /* control_fsm_rtl.vhd:192:50  */
  assign n2704_o = s_command == 8'b01010100;
  /* control_fsm_rtl.vhd:191:67  */
  assign n2705_o = n2704_o ? 7'b0001101 : n2709_o;
  /* control_fsm_rtl.vhd:193:50  */
  assign n2708_o = s_command == 8'b01010010;
  /* control_fsm_rtl.vhd:192:67  */
  assign n2709_o = n2708_o ? 7'b0001110 : n2713_o;
  /* control_fsm_rtl.vhd:194:50  */
  assign n2712_o = s_command == 8'b01010011;
  /* control_fsm_rtl.vhd:193:67  */
  assign n2713_o = n2712_o ? 7'b0001111 : n2717_o;
  /* control_fsm_rtl.vhd:195:50  */
  assign n2716_o = s_command == 8'b10000010;
  /* control_fsm_rtl.vhd:194:67  */
  assign n2717_o = n2716_o ? 7'b0010000 : n2721_o;
  /* control_fsm_rtl.vhd:196:50  */
  assign n2720_o = s_command == 8'b10110000;
  /* control_fsm_rtl.vhd:195:67  */
  assign n2721_o = n2720_o ? 7'b0010001 : n2725_o;
  /* control_fsm_rtl.vhd:197:50  */
  assign n2724_o = s_command == 8'b10110101;
  /* control_fsm_rtl.vhd:196:67  */
  assign n2725_o = n2724_o ? 7'b0010010 : n2729_o;
  /* control_fsm_rtl.vhd:198:50  */
  assign n2728_o = s_command == 8'b10110100;
  /* control_fsm_rtl.vhd:197:67  */
  assign n2729_o = n2728_o ? 7'b0010011 : n2734_o;
  /* control_fsm_rtl.vhd:199:37  */
  assign n2731_o = s_command[7:3];
  /* control_fsm_rtl.vhd:199:50  */
  assign n2733_o = n2731_o == 5'b10111;
  /* control_fsm_rtl.vhd:198:67  */
  assign n2734_o = n2733_o ? 7'b0010100 : n2739_o;
  /* control_fsm_rtl.vhd:200:37  */
  assign n2736_o = s_command[7:1];
  /* control_fsm_rtl.vhd:200:50  */
  assign n2738_o = n2736_o == 7'b1011011;
  /* control_fsm_rtl.vhd:199:67  */
  assign n2739_o = n2738_o ? 7'b0010101 : n2743_o;
  /* control_fsm_rtl.vhd:201:50  */
  assign n2742_o = s_command == 8'b11100100;
  /* control_fsm_rtl.vhd:200:67  */
  assign n2743_o = n2742_o ? 7'b0010110 : n2747_o;
  /* control_fsm_rtl.vhd:202:50  */
  assign n2746_o = s_command == 8'b11000011;
  /* control_fsm_rtl.vhd:201:67  */
  assign n2747_o = n2746_o ? 7'b0010111 : n2751_o;
  /* control_fsm_rtl.vhd:203:50  */
  assign n2750_o = s_command == 8'b11000010;
  /* control_fsm_rtl.vhd:202:67  */
  assign n2751_o = n2750_o ? 7'b0011000 : n2755_o;
  /* control_fsm_rtl.vhd:204:50  */
  assign n2754_o = s_command == 8'b11110100;
  /* control_fsm_rtl.vhd:203:67  */
  assign n2755_o = n2754_o ? 7'b0011001 : n2759_o;
  /* control_fsm_rtl.vhd:205:50  */
  assign n2758_o = s_command == 8'b10110011;
  /* control_fsm_rtl.vhd:204:67  */
  assign n2759_o = n2758_o ? 7'b0011010 : n2763_o;
  /* control_fsm_rtl.vhd:206:50  */
  assign n2762_o = s_command == 8'b10110010;
  /* control_fsm_rtl.vhd:205:67  */
  assign n2763_o = n2762_o ? 7'b0011011 : n2767_o;
  /* control_fsm_rtl.vhd:207:50  */
  assign n2766_o = s_command == 8'b11010100;
  /* control_fsm_rtl.vhd:206:67  */
  assign n2767_o = n2766_o ? 7'b0011100 : n2771_o;
  /* control_fsm_rtl.vhd:208:50  */
  assign n2770_o = s_command == 8'b00010100;
  /* control_fsm_rtl.vhd:207:67  */
  assign n2771_o = n2770_o ? 7'b0011101 : n2776_o;
  /* control_fsm_rtl.vhd:209:37  */
  assign n2773_o = s_command[7:3];
  /* control_fsm_rtl.vhd:209:50  */
  assign n2775_o = n2773_o == 5'b00011;
  /* control_fsm_rtl.vhd:208:67  */
  assign n2776_o = n2775_o ? 7'b0011110 : n2780_o;
  /* control_fsm_rtl.vhd:210:50  */
  assign n2779_o = s_command == 8'b00010101;
  /* control_fsm_rtl.vhd:209:67  */
  assign n2780_o = n2779_o ? 7'b0011111 : n2785_o;
  /* control_fsm_rtl.vhd:211:37  */
  assign n2782_o = s_command[7:1];
  /* control_fsm_rtl.vhd:211:50  */
  assign n2784_o = n2782_o == 7'b0001011;
  /* control_fsm_rtl.vhd:210:67  */
  assign n2785_o = n2784_o ? 7'b0100000 : n2789_o;
  /* control_fsm_rtl.vhd:212:50  */
  assign n2788_o = s_command == 8'b10000100;
  /* control_fsm_rtl.vhd:211:67  */
  assign n2789_o = n2788_o ? 7'b0100001 : n2794_o;
  /* control_fsm_rtl.vhd:213:37  */
  assign n2791_o = s_command[7:3];
  /* control_fsm_rtl.vhd:213:50  */
  assign n2793_o = n2791_o == 5'b11011;
  /* control_fsm_rtl.vhd:212:67  */
  assign n2794_o = n2793_o ? 7'b0100010 : n2798_o;
  /* control_fsm_rtl.vhd:214:50  */
  assign n2797_o = s_command == 8'b11010101;
  /* control_fsm_rtl.vhd:213:67  */
  assign n2798_o = n2797_o ? 7'b0100011 : n2802_o;
  /* control_fsm_rtl.vhd:215:50  */
  assign n2801_o = s_command == 8'b00000100;
  /* control_fsm_rtl.vhd:214:67  */
  assign n2802_o = n2801_o ? 7'b0100100 : n2807_o;
  /* control_fsm_rtl.vhd:216:37  */
  assign n2804_o = s_command[7:3];
  /* control_fsm_rtl.vhd:216:50  */
  assign n2806_o = n2804_o == 5'b00001;
  /* control_fsm_rtl.vhd:215:67  */
  assign n2807_o = n2806_o ? 7'b0100101 : n2811_o;
  /* control_fsm_rtl.vhd:217:50  */
  assign n2810_o = s_command == 8'b00000101;
  /* control_fsm_rtl.vhd:216:67  */
  assign n2811_o = n2810_o ? 7'b0100110 : n2816_o;
  /* control_fsm_rtl.vhd:218:37  */
  assign n2813_o = s_command[7:1];
  /* control_fsm_rtl.vhd:218:50  */
  assign n2815_o = n2813_o == 7'b0000011;
  /* control_fsm_rtl.vhd:217:67  */
  assign n2816_o = n2815_o ? 7'b0100111 : n2820_o;
  /* control_fsm_rtl.vhd:219:50  */
  assign n2819_o = s_command == 8'b10100011;
  /* control_fsm_rtl.vhd:218:67  */
  assign n2820_o = n2819_o ? 7'b0101000 : n2824_o;
  /* control_fsm_rtl.vhd:220:50  */
  assign n2823_o = s_command == 8'b00100000;
  /* control_fsm_rtl.vhd:219:67  */
  assign n2824_o = n2823_o ? 7'b0101001 : n2828_o;
  /* control_fsm_rtl.vhd:221:50  */
  assign n2827_o = s_command == 8'b00010000;
  /* control_fsm_rtl.vhd:220:67  */
  assign n2828_o = n2827_o ? 7'b0101010 : n2832_o;
  /* control_fsm_rtl.vhd:222:50  */
  assign n2831_o = s_command == 8'b01000000;
  /* control_fsm_rtl.vhd:221:67  */
  assign n2832_o = n2831_o ? 7'b0101011 : n2836_o;
  /* control_fsm_rtl.vhd:223:50  */
  assign n2835_o = s_command == 8'b01110011;
  /* control_fsm_rtl.vhd:222:67  */
  assign n2836_o = n2835_o ? 7'b0101100 : n2840_o;
  /* control_fsm_rtl.vhd:224:50  */
  assign n2839_o = s_command == 8'b00110000;
  /* control_fsm_rtl.vhd:223:67  */
  assign n2840_o = n2839_o ? 7'b0101101 : n2844_o;
  /* control_fsm_rtl.vhd:225:50  */
  assign n2843_o = s_command == 8'b01010000;
  /* control_fsm_rtl.vhd:224:67  */
  assign n2844_o = n2843_o ? 7'b0101110 : n2848_o;
  /* control_fsm_rtl.vhd:226:50  */
  assign n2847_o = s_command == 8'b01110000;
  /* control_fsm_rtl.vhd:225:67  */
  assign n2848_o = n2847_o ? 7'b0101111 : n2852_o;
  /* control_fsm_rtl.vhd:227:50  */
  assign n2851_o = s_command == 8'b01100000;
  /* control_fsm_rtl.vhd:226:67  */
  assign n2852_o = n2851_o ? 7'b0110000 : n2856_o;
  /* control_fsm_rtl.vhd:228:50  */
  assign n2855_o = s_command == 8'b00010010;
  /* control_fsm_rtl.vhd:227:67  */
  assign n2856_o = n2855_o ? 7'b0110001 : n2860_o;
  /* control_fsm_rtl.vhd:229:50  */
  assign n2859_o = s_command == 8'b00000010;
  /* control_fsm_rtl.vhd:228:67  */
  assign n2860_o = n2859_o ? 7'b0110010 : n2865_o;
  /* control_fsm_rtl.vhd:230:37  */
  assign n2862_o = s_command[7:3];
  /* control_fsm_rtl.vhd:230:50  */
  assign n2864_o = n2862_o == 5'b11101;
  /* control_fsm_rtl.vhd:229:67  */
  assign n2865_o = n2864_o ? 7'b0110011 : n2869_o;
  /* control_fsm_rtl.vhd:231:50  */
  assign n2868_o = s_command == 8'b11100101;
  /* control_fsm_rtl.vhd:230:67  */
  assign n2869_o = n2868_o ? 7'b0110100 : n2874_o;
  /* control_fsm_rtl.vhd:232:37  */
  assign n2871_o = s_command[7:1];
  /* control_fsm_rtl.vhd:232:50  */
  assign n2873_o = n2871_o == 7'b1110011;
  /* control_fsm_rtl.vhd:231:67  */
  assign n2874_o = n2873_o ? 7'b0110101 : n2878_o;
  /* control_fsm_rtl.vhd:233:50  */
  assign n2877_o = s_command == 8'b01110100;
  /* control_fsm_rtl.vhd:232:67  */
  assign n2878_o = n2877_o ? 7'b0110110 : n2883_o;
  /* control_fsm_rtl.vhd:234:37  */
  assign n2880_o = s_command[7:3];
  /* control_fsm_rtl.vhd:234:50  */
  assign n2882_o = n2880_o == 5'b11111;
  /* control_fsm_rtl.vhd:233:67  */
  assign n2883_o = n2882_o ? 7'b0110111 : n2888_o;
  /* control_fsm_rtl.vhd:235:37  */
  assign n2885_o = s_command[7:3];
  /* control_fsm_rtl.vhd:235:50  */
  assign n2887_o = n2885_o == 5'b10101;
  /* control_fsm_rtl.vhd:234:67  */
  assign n2888_o = n2887_o ? 7'b0111000 : n2893_o;
  /* control_fsm_rtl.vhd:236:37  */
  assign n2890_o = s_command[7:3];
  /* control_fsm_rtl.vhd:236:50  */
  assign n2892_o = n2890_o == 5'b01111;
  /* control_fsm_rtl.vhd:235:67  */
  assign n2893_o = n2892_o ? 7'b0111001 : n2897_o;
  /* control_fsm_rtl.vhd:237:50  */
  assign n2896_o = s_command == 8'b11110101;
  /* control_fsm_rtl.vhd:236:67  */
  assign n2897_o = n2896_o ? 7'b0111010 : n2902_o;
  /* control_fsm_rtl.vhd:238:37  */
  assign n2899_o = s_command[7:3];
  /* control_fsm_rtl.vhd:238:50  */
  assign n2901_o = n2899_o == 5'b10001;
  /* control_fsm_rtl.vhd:237:67  */
  assign n2902_o = n2901_o ? 7'b0111011 : n2906_o;
  /* control_fsm_rtl.vhd:239:50  */
  assign n2905_o = s_command == 8'b10000101;
  /* control_fsm_rtl.vhd:238:67  */
  assign n2906_o = n2905_o ? 7'b0111100 : n2911_o;
  /* control_fsm_rtl.vhd:240:37  */
  assign n2908_o = s_command[7:1];
  /* control_fsm_rtl.vhd:240:50  */
  assign n2910_o = n2908_o == 7'b1000011;
  /* control_fsm_rtl.vhd:239:67  */
  assign n2911_o = n2910_o ? 7'b0111101 : n2915_o;
  /* control_fsm_rtl.vhd:241:50  */
  assign n2914_o = s_command == 8'b01110101;
  /* control_fsm_rtl.vhd:240:67  */
  assign n2915_o = n2914_o ? 7'b0111110 : n2920_o;
  /* control_fsm_rtl.vhd:242:37  */
  assign n2917_o = s_command[7:1];
  /* control_fsm_rtl.vhd:242:50  */
  assign n2919_o = n2917_o == 7'b1111011;
  /* control_fsm_rtl.vhd:241:67  */
  assign n2920_o = n2919_o ? 7'b0111111 : n2925_o;
  /* control_fsm_rtl.vhd:243:37  */
  assign n2922_o = s_command[7:1];
  /* control_fsm_rtl.vhd:243:50  */
  assign n2924_o = n2922_o == 7'b1010011;
  /* control_fsm_rtl.vhd:242:67  */
  assign n2925_o = n2924_o ? 7'b1000000 : n2930_o;
  /* control_fsm_rtl.vhd:244:37  */
  assign n2927_o = s_command[7:1];
  /* control_fsm_rtl.vhd:244:50  */
  assign n2929_o = n2927_o == 7'b0111011;
  /* control_fsm_rtl.vhd:243:67  */
  assign n2930_o = n2929_o ? 7'b1000001 : n2934_o;
  /* control_fsm_rtl.vhd:245:50  */
  assign n2933_o = s_command == 8'b10010011;
  /* control_fsm_rtl.vhd:244:67  */
  assign n2934_o = n2933_o ? 7'b1000010 : n2938_o;
  /* control_fsm_rtl.vhd:246:50  */
  assign n2937_o = s_command == 8'b10000011;
  /* control_fsm_rtl.vhd:245:67  */
  assign n2938_o = n2937_o ? 7'b1000011 : n2943_o;
  /* control_fsm_rtl.vhd:247:37  */
  assign n2940_o = s_command[7:1];
  /* control_fsm_rtl.vhd:247:50  */
  assign n2942_o = n2940_o == 7'b1110001;
  /* control_fsm_rtl.vhd:246:67  */
  assign n2943_o = n2942_o ? 7'b1000100 : n2947_o;
  /* control_fsm_rtl.vhd:248:50  */
  assign n2946_o = s_command == 8'b11100000;
  /* control_fsm_rtl.vhd:247:67  */
  assign n2947_o = n2946_o ? 7'b1000101 : n2952_o;
  /* control_fsm_rtl.vhd:249:37  */
  assign n2949_o = s_command[7:1];
  /* control_fsm_rtl.vhd:249:50  */
  assign n2951_o = n2949_o == 7'b1111001;
  /* control_fsm_rtl.vhd:248:67  */
  assign n2952_o = n2951_o ? 7'b1000110 : n2956_o;
  /* control_fsm_rtl.vhd:250:50  */
  assign n2955_o = s_command == 8'b11110000;
  /* control_fsm_rtl.vhd:249:67  */
  assign n2956_o = n2955_o ? 7'b1000111 : n2960_o;
  /* control_fsm_rtl.vhd:251:50  */
  assign n2959_o = s_command == 8'b10100010;
  /* control_fsm_rtl.vhd:250:67  */
  assign n2960_o = n2959_o ? 7'b1001000 : n2964_o;
  /* control_fsm_rtl.vhd:252:50  */
  assign n2963_o = s_command == 8'b10010010;
  /* control_fsm_rtl.vhd:251:67  */
  assign n2964_o = n2963_o ? 7'b1001001 : n2968_o;
  /* control_fsm_rtl.vhd:253:50  */
  assign n2967_o = s_command == 8'b10010000;
  /* control_fsm_rtl.vhd:252:67  */
  assign n2968_o = n2967_o ? 7'b1001010 : n2972_o;
  /* control_fsm_rtl.vhd:254:50  */
  assign n2971_o = s_command == 8'b10100100;
  /* control_fsm_rtl.vhd:253:67  */
  assign n2972_o = n2971_o ? 7'b1001011 : n2976_o;
  /* control_fsm_rtl.vhd:255:50  */
  assign n2975_o = s_command == 8'b00000000;
  /* control_fsm_rtl.vhd:254:67  */
  assign n2976_o = n2975_o ? 7'b1001100 : n2981_o;
  /* control_fsm_rtl.vhd:256:37  */
  assign n2978_o = s_command[7:3];
  /* control_fsm_rtl.vhd:256:50  */
  assign n2980_o = n2978_o == 5'b01001;
  /* control_fsm_rtl.vhd:255:67  */
  assign n2981_o = n2980_o ? 7'b1001101 : n2985_o;
  /* control_fsm_rtl.vhd:257:50  */
  assign n2984_o = s_command == 8'b01000101;
  /* control_fsm_rtl.vhd:256:67  */
  assign n2985_o = n2984_o ? 7'b1001110 : n2990_o;
  /* control_fsm_rtl.vhd:258:37  */
  assign n2987_o = s_command[7:1];
  /* control_fsm_rtl.vhd:258:50  */
  assign n2989_o = n2987_o == 7'b0100011;
  /* control_fsm_rtl.vhd:257:67  */
  assign n2990_o = n2989_o ? 7'b1001111 : n2994_o;
  /* control_fsm_rtl.vhd:259:50  */
  assign n2993_o = s_command == 8'b01000100;
  /* control_fsm_rtl.vhd:258:67  */
  assign n2994_o = n2993_o ? 7'b1010000 : n2998_o;
  /* control_fsm_rtl.vhd:260:50  */
  assign n2997_o = s_command == 8'b01000010;
  /* control_fsm_rtl.vhd:259:67  */
  assign n2998_o = n2997_o ? 7'b1010001 : n3002_o;
  /* control_fsm_rtl.vhd:261:50  */
  assign n3001_o = s_command == 8'b01000011;
  /* control_fsm_rtl.vhd:260:67  */
  assign n3002_o = n3001_o ? 7'b1010010 : n3006_o;
  /* control_fsm_rtl.vhd:262:50  */
  assign n3005_o = s_command == 8'b01110010;
  /* control_fsm_rtl.vhd:261:67  */
  assign n3006_o = n3005_o ? 7'b1010011 : n3010_o;
  /* control_fsm_rtl.vhd:263:50  */
  assign n3009_o = s_command == 8'b10100000;
  /* control_fsm_rtl.vhd:262:67  */
  assign n3010_o = n3009_o ? 7'b1010100 : n3014_o;
  /* control_fsm_rtl.vhd:264:50  */
  assign n3013_o = s_command == 8'b11010000;
  /* control_fsm_rtl.vhd:263:67  */
  assign n3014_o = n3013_o ? 7'b1010101 : n3018_o;
  /* control_fsm_rtl.vhd:265:50  */
  assign n3017_o = s_command == 8'b11000000;
  /* control_fsm_rtl.vhd:264:67  */
  assign n3018_o = n3017_o ? 7'b1010110 : n3022_o;
  /* control_fsm_rtl.vhd:266:50  */
  assign n3021_o = s_command == 8'b00100010;
  /* control_fsm_rtl.vhd:265:67  */
  assign n3022_o = n3021_o ? 7'b1010111 : n3026_o;
  /* control_fsm_rtl.vhd:267:50  */
  assign n3025_o = s_command == 8'b00110010;
  /* control_fsm_rtl.vhd:266:67  */
  assign n3026_o = n3025_o ? 7'b1011000 : n3030_o;
  /* control_fsm_rtl.vhd:268:50  */
  assign n3029_o = s_command == 8'b00100011;
  /* control_fsm_rtl.vhd:267:67  */
  assign n3030_o = n3029_o ? 7'b1011001 : n3034_o;
  /* control_fsm_rtl.vhd:269:50  */
  assign n3033_o = s_command == 8'b00110011;
  /* control_fsm_rtl.vhd:268:67  */
  assign n3034_o = n3033_o ? 7'b1011010 : n3038_o;
  /* control_fsm_rtl.vhd:270:50  */
  assign n3037_o = s_command == 8'b00000011;
  /* control_fsm_rtl.vhd:269:67  */
  assign n3038_o = n3037_o ? 7'b1011011 : n3042_o;
  /* control_fsm_rtl.vhd:271:50  */
  assign n3041_o = s_command == 8'b00010011;
  /* control_fsm_rtl.vhd:270:67  */
  assign n3042_o = n3041_o ? 7'b1011100 : n3046_o;
  /* control_fsm_rtl.vhd:272:50  */
  assign n3045_o = s_command == 8'b11010011;
  /* control_fsm_rtl.vhd:271:67  */
  assign n3046_o = n3045_o ? 7'b1011101 : n3050_o;
  /* control_fsm_rtl.vhd:273:50  */
  assign n3049_o = s_command == 8'b11010010;
  /* control_fsm_rtl.vhd:272:67  */
  assign n3050_o = n3049_o ? 7'b1011110 : n3054_o;
  /* control_fsm_rtl.vhd:274:50  */
  assign n3053_o = s_command == 8'b10000000;
  /* control_fsm_rtl.vhd:273:67  */
  assign n3054_o = n3053_o ? 7'b1011111 : n3059_o;
  /* control_fsm_rtl.vhd:275:37  */
  assign n3056_o = s_command[7:3];
  /* control_fsm_rtl.vhd:275:50  */
  assign n3058_o = n3056_o == 5'b10011;
  /* control_fsm_rtl.vhd:274:67  */
  assign n3059_o = n3058_o ? 7'b1100000 : n3063_o;
  /* control_fsm_rtl.vhd:276:50  */
  assign n3062_o = s_command == 8'b10010101;
  /* control_fsm_rtl.vhd:275:67  */
  assign n3063_o = n3062_o ? 7'b1100001 : n3068_o;
  /* control_fsm_rtl.vhd:277:37  */
  assign n3065_o = s_command[7:1];
  /* control_fsm_rtl.vhd:277:50  */
  assign n3067_o = n3065_o == 7'b1001011;
  /* control_fsm_rtl.vhd:276:67  */
  assign n3068_o = n3067_o ? 7'b1100010 : n3072_o;
  /* control_fsm_rtl.vhd:278:50  */
  assign n3071_o = s_command == 8'b10010100;
  /* control_fsm_rtl.vhd:277:67  */
  assign n3072_o = n3071_o ? 7'b1100011 : n3076_o;
  /* control_fsm_rtl.vhd:279:50  */
  assign n3075_o = s_command == 8'b11000100;
  /* control_fsm_rtl.vhd:278:67  */
  assign n3076_o = n3075_o ? 7'b1100100 : n3081_o;
  /* control_fsm_rtl.vhd:280:37  */
  assign n3078_o = s_command[7:3];
  /* control_fsm_rtl.vhd:280:50  */
  assign n3080_o = n3078_o == 5'b11001;
  /* control_fsm_rtl.vhd:279:67  */
  assign n3081_o = n3080_o ? 7'b1100101 : n3085_o;
  /* control_fsm_rtl.vhd:281:50  */
  assign n3084_o = s_command == 8'b11000101;
  /* control_fsm_rtl.vhd:280:67  */
  assign n3085_o = n3084_o ? 7'b1100110 : n3090_o;
  /* control_fsm_rtl.vhd:282:37  */
  assign n3087_o = s_command[7:1];
  /* control_fsm_rtl.vhd:282:50  */
  assign n3089_o = n3087_o == 7'b1100011;
  /* control_fsm_rtl.vhd:281:67  */
  assign n3090_o = n3089_o ? 7'b1100111 : n3095_o;
  /* control_fsm_rtl.vhd:283:37  */
  assign n3092_o = s_command[7:1];
  /* control_fsm_rtl.vhd:283:50  */
  assign n3094_o = n3092_o == 7'b1101011;
  /* control_fsm_rtl.vhd:282:67  */
  assign n3095_o = n3094_o ? 7'b1101000 : n3100_o;
  /* control_fsm_rtl.vhd:284:37  */
  assign n3097_o = s_command[7:3];
  /* control_fsm_rtl.vhd:284:50  */
  assign n3099_o = n3097_o == 5'b01101;
  /* control_fsm_rtl.vhd:283:67  */
  assign n3100_o = n3099_o ? 7'b1101001 : n3104_o;
  /* control_fsm_rtl.vhd:285:50  */
  assign n3103_o = s_command == 8'b01100101;
  /* control_fsm_rtl.vhd:284:67  */
  assign n3104_o = n3103_o ? 7'b1101010 : n3109_o;
  /* control_fsm_rtl.vhd:286:37  */
  assign n3106_o = s_command[7:1];
  /* control_fsm_rtl.vhd:286:50  */
  assign n3108_o = n3106_o == 7'b0110011;
  /* control_fsm_rtl.vhd:285:67  */
  assign n3109_o = n3108_o ? 7'b1101011 : n3113_o;
  /* control_fsm_rtl.vhd:287:50  */
  assign n3112_o = s_command == 8'b01100100;
  /* control_fsm_rtl.vhd:286:67  */
  assign n3113_o = n3112_o ? 7'b1101100 : n3117_o;
  /* control_fsm_rtl.vhd:288:50  */
  assign n3116_o = s_command == 8'b01100010;
  /* control_fsm_rtl.vhd:287:67  */
  assign n3117_o = n3116_o ? 7'b1101101 : n3121_o;
  /* control_fsm_rtl.vhd:289:50  */
  assign n3120_o = s_command == 8'b01100011;
  /* control_fsm_rtl.vhd:288:67  */
  assign n3121_o = n3120_o ? 7'b1101110 : 7'b1001100;
  /* control_fsm_rtl.vhd:334:13  */
  assign n3125_o = state == 3'b000;
  /* control_fsm_rtl.vhd:340:21  */
  assign n3126_o = ~intblock_i;
  /* control_fsm_rtl.vhd:340:48  */
  assign n3128_o = s_instr_category != 7'b1011000;
  /* control_fsm_rtl.vhd:340:27  */
  assign n3129_o = n3126_o & n3128_o;
  /* control_fsm_rtl.vhd:343:34  */
  assign n3131_o = state == 3'b001;
  /* control_fsm_rtl.vhd:343:25  */
  assign n3132_o = s_intpre & n3131_o;
  /* control_fsm_rtl.vhd:343:42  */
  assign n3133_o = n3132_o | s_intpre2;
  /* control_fsm_rtl.vhd:340:59  */
  assign n3134_o = n3129_o & n3133_o;
  /* control_fsm_rtl.vhd:344:17  */
  assign n3136_o = state == 3'b001;
  /* control_fsm_rtl.vhd:349:20  */
  assign n3138_o = state == 3'b010;
  /* control_fsm_rtl.vhd:350:19  */
  assign n3139_o = n2641_o & n2636_o;
  /* control_fsm_rtl.vhd:350:27  */
  assign n3140_o = n3139_o & s_ie0;
  /* control_fsm_rtl.vhd:358:22  */
  assign n3141_o = n2640_o & n2635_o;
  /* control_fsm_rtl.vhd:358:30  */
  assign n3142_o = n3141_o & s_tf0;
  /* control_fsm_rtl.vhd:364:22  */
  assign n3143_o = n2639_o & n2634_o;
  /* control_fsm_rtl.vhd:364:30  */
  assign n3144_o = n3143_o & s_ie1;
  /* control_fsm_rtl.vhd:372:22  */
  assign n3145_o = n2638_o & n2633_o;
  /* control_fsm_rtl.vhd:372:30  */
  assign n3146_o = n3145_o & s_tf1;
  /* control_fsm_rtl.vhd:378:22  */
  assign n3147_o = n2637_o & n2632_o;
  /* control_fsm_rtl.vhd:378:39  */
  assign n3148_o = s_ri | s_ti;
  /* control_fsm_rtl.vhd:378:29  */
  assign n3149_o = n3147_o & n3148_o;
  /* control_fsm_rtl.vhd:382:21  */
  assign n3150_o = n2636_o & s_ie0;
  /* control_fsm_rtl.vhd:390:22  */
  assign n3151_o = n2635_o & s_tf0;
  /* control_fsm_rtl.vhd:396:22  */
  assign n3152_o = n2634_o & s_ie1;
  /* control_fsm_rtl.vhd:404:22  */
  assign n3153_o = n2633_o & s_tf1;
  /* control_fsm_rtl.vhd:410:31  */
  assign n3154_o = s_ri | s_ti;
  /* control_fsm_rtl.vhd:410:21  */
  assign n3155_o = n2632_o & n3154_o;
  /* control_fsm_rtl.vhd:410:11  */
  assign n3158_o = n3155_o ? 4'b1001 : 4'b0000;
  /* control_fsm_rtl.vhd:410:11  */
  assign n3161_o = n3155_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:410:11  */
  assign n3164_o = n3155_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:404:11  */
  assign n3167_o = n3153_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:404:11  */
  assign n3170_o = n3153_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:404:11  */
  assign n3172_o = n3153_o ? 4'b1000 : n3158_o;
  /* control_fsm_rtl.vhd:404:11  */
  assign n3174_o = n3153_o ? 1'b1 : n3161_o;
  /* control_fsm_rtl.vhd:404:11  */
  assign n3176_o = n3153_o ? 1'b1 : n3164_o;
  /* control_fsm_rtl.vhd:396:11  */
  assign n3178_o = n3152_o ? 3'b110 : n3167_o;
  /* control_fsm_rtl.vhd:396:11  */
  assign n3180_o = n3152_o ? 4'b0011 : n3170_o;
  /* control_fsm_rtl.vhd:396:11  */
  assign n3182_o = n3152_o ? 4'b0111 : n3172_o;
  /* control_fsm_rtl.vhd:396:11  */
  assign n3184_o = n3152_o ? 1'b1 : n3174_o;
  /* control_fsm_rtl.vhd:396:11  */
  assign n3186_o = n3152_o ? 1'b1 : n3176_o;
  /* control_fsm_rtl.vhd:396:11  */
  assign n3189_o = n3152_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:396:11  */
  assign n3192_o = n3152_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:390:11  */
  assign n3194_o = n3151_o ? 3'b110 : n3178_o;
  /* control_fsm_rtl.vhd:390:11  */
  assign n3196_o = n3151_o ? 4'b0010 : n3180_o;
  /* control_fsm_rtl.vhd:390:11  */
  assign n3198_o = n3151_o ? 4'b0110 : n3182_o;
  /* control_fsm_rtl.vhd:390:11  */
  assign n3200_o = n3151_o ? 1'b1 : n3184_o;
  /* control_fsm_rtl.vhd:390:11  */
  assign n3202_o = n3151_o ? 1'b1 : n3186_o;
  /* control_fsm_rtl.vhd:390:11  */
  assign n3204_o = n3151_o ? 1'b0 : n3189_o;
  /* control_fsm_rtl.vhd:390:11  */
  assign n3206_o = n3151_o ? 1'b0 : n3192_o;
  /* control_fsm_rtl.vhd:382:10  */
  assign n3208_o = n3150_o ? 3'b110 : n3194_o;
  /* control_fsm_rtl.vhd:382:10  */
  assign n3210_o = n3150_o ? 4'b0001 : n3196_o;
  /* control_fsm_rtl.vhd:382:10  */
  assign n3212_o = n3150_o ? 4'b0101 : n3198_o;
  /* control_fsm_rtl.vhd:382:10  */
  assign n3214_o = n3150_o ? 1'b1 : n3200_o;
  /* control_fsm_rtl.vhd:382:10  */
  assign n3216_o = n3150_o ? 1'b1 : n3202_o;
  /* control_fsm_rtl.vhd:382:10  */
  assign n3219_o = n3150_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:382:10  */
  assign n3221_o = n3150_o ? 1'b0 : n3204_o;
  /* control_fsm_rtl.vhd:382:10  */
  assign n3224_o = n3150_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:382:10  */
  assign n3226_o = n3150_o ? 1'b0 : n3206_o;
  /* control_fsm_rtl.vhd:378:11  */
  assign n3228_o = n3149_o ? 3'b000 : n3208_o;
  /* control_fsm_rtl.vhd:378:11  */
  assign n3230_o = n3149_o ? 4'b0000 : n3210_o;
  /* control_fsm_rtl.vhd:378:11  */
  assign n3232_o = n3149_o ? 4'b1001 : n3212_o;
  /* control_fsm_rtl.vhd:378:11  */
  assign n3234_o = n3149_o ? 1'b0 : n3214_o;
  /* control_fsm_rtl.vhd:378:11  */
  assign n3236_o = n3149_o ? 1'b0 : n3216_o;
  /* control_fsm_rtl.vhd:378:11  */
  assign n3239_o = n3149_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:378:11  */
  assign n3242_o = n3149_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:378:11  */
  assign n3244_o = n3149_o ? 1'b0 : n3219_o;
  /* control_fsm_rtl.vhd:378:11  */
  assign n3246_o = n3149_o ? 1'b0 : n3221_o;
  /* control_fsm_rtl.vhd:378:11  */
  assign n3248_o = n3149_o ? 1'b0 : n3224_o;
  /* control_fsm_rtl.vhd:378:11  */
  assign n3250_o = n3149_o ? 1'b0 : n3226_o;
  /* control_fsm_rtl.vhd:372:11  */
  assign n3252_o = n3146_o ? 3'b110 : n3228_o;
  /* control_fsm_rtl.vhd:372:11  */
  assign n3254_o = n3146_o ? 4'b0100 : n3230_o;
  /* control_fsm_rtl.vhd:372:11  */
  assign n3256_o = n3146_o ? 4'b1000 : n3232_o;
  /* control_fsm_rtl.vhd:372:11  */
  assign n3258_o = n3146_o ? 1'b0 : n3234_o;
  /* control_fsm_rtl.vhd:372:11  */
  assign n3260_o = n3146_o ? 1'b0 : n3236_o;
  /* control_fsm_rtl.vhd:372:11  */
  assign n3262_o = n3146_o ? 1'b1 : n3239_o;
  /* control_fsm_rtl.vhd:372:11  */
  assign n3264_o = n3146_o ? 1'b1 : n3242_o;
  /* control_fsm_rtl.vhd:372:11  */
  assign n3266_o = n3146_o ? 1'b0 : n3244_o;
  /* control_fsm_rtl.vhd:372:11  */
  assign n3268_o = n3146_o ? 1'b0 : n3246_o;
  /* control_fsm_rtl.vhd:372:11  */
  assign n3270_o = n3146_o ? 1'b0 : n3248_o;
  /* control_fsm_rtl.vhd:372:11  */
  assign n3272_o = n3146_o ? 1'b0 : n3250_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3274_o = n3144_o ? 3'b110 : n3252_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3276_o = n3144_o ? 4'b0011 : n3254_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3278_o = n3144_o ? 4'b0111 : n3256_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3280_o = n3144_o ? 1'b0 : n3258_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3282_o = n3144_o ? 1'b0 : n3260_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3284_o = n3144_o ? 1'b1 : n3262_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3286_o = n3144_o ? 1'b1 : n3264_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3288_o = n3144_o ? 1'b0 : n3266_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3290_o = n3144_o ? 1'b0 : n3268_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3293_o = n3144_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3295_o = n3144_o ? 1'b0 : n3270_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3297_o = n3144_o ? 1'b0 : n3272_o;
  /* control_fsm_rtl.vhd:364:11  */
  assign n3300_o = n3144_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3302_o = n3142_o ? 3'b110 : n3274_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3304_o = n3142_o ? 4'b0010 : n3276_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3306_o = n3142_o ? 4'b0110 : n3278_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3308_o = n3142_o ? 1'b0 : n3280_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3310_o = n3142_o ? 1'b0 : n3282_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3312_o = n3142_o ? 1'b1 : n3284_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3314_o = n3142_o ? 1'b1 : n3286_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3316_o = n3142_o ? 1'b0 : n3288_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3318_o = n3142_o ? 1'b0 : n3290_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3320_o = n3142_o ? 1'b0 : n3293_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3322_o = n3142_o ? 1'b0 : n3295_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3324_o = n3142_o ? 1'b0 : n3297_o;
  /* control_fsm_rtl.vhd:358:11  */
  assign n3326_o = n3142_o ? 1'b0 : n3300_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3328_o = n3140_o ? 3'b110 : n3302_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3330_o = n3140_o ? 4'b0001 : n3304_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3332_o = n3140_o ? 4'b0101 : n3306_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3334_o = n3140_o ? 1'b0 : n3308_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3336_o = n3140_o ? 1'b0 : n3310_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3338_o = n3140_o ? 1'b1 : n3312_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3340_o = n3140_o ? 1'b1 : n3314_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3342_o = n3140_o ? 1'b0 : n3316_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3344_o = n3140_o ? 1'b0 : n3318_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3347_o = n3140_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3349_o = n3140_o ? 1'b0 : n3320_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3351_o = n3140_o ? 1'b0 : n3322_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3353_o = n3140_o ? 1'b0 : n3324_o;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3356_o = n3140_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:350:11  */
  assign n3358_o = n3140_o ? 1'b0 : n3326_o;
  /* control_fsm_rtl.vhd:418:20  */
  assign n3360_o = state == 3'b011;
  /* control_fsm_rtl.vhd:423:20  */
  assign n3362_o = state == 3'b100;
  /* control_fsm_rtl.vhd:423:9  */
  assign n3365_o = n3362_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:423:9  */
  assign n3368_o = n3362_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:423:9  */
  assign n3371_o = n3362_o ? 4'b0010 : 4'b0000;
  /* control_fsm_rtl.vhd:423:9  */
  assign n3374_o = n3362_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:423:9  */
  assign n3377_o = n3362_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:418:9  */
  assign n3380_o = n3360_o ? 3'b100 : 3'b001;
  /* control_fsm_rtl.vhd:418:9  */
  assign n3382_o = n3360_o ? 4'b0000 : n3365_o;
  /* control_fsm_rtl.vhd:418:9  */
  assign n3384_o = n3360_o ? 3'b101 : n3368_o;
  /* control_fsm_rtl.vhd:418:9  */
  assign n3386_o = n3360_o ? 4'b0001 : n3371_o;
  /* control_fsm_rtl.vhd:418:9  */
  assign n3388_o = n3360_o ? 4'b0101 : n3374_o;
  /* control_fsm_rtl.vhd:418:9  */
  assign n3390_o = n3360_o ? 1'b0 : n3377_o;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3392_o = n3138_o ? 3'b011 : n3380_o;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3394_o = n3138_o ? 4'b0000 : n3382_o;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3395_o = n3138_o ? n3328_o : n3384_o;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3397_o = n3138_o ? 4'b0000 : n3386_o;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3398_o = n3138_o ? n3330_o : n3388_o;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3400_o = n3138_o ? n3332_o : 4'b0000;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3402_o = n3138_o ? 1'b0 : n3390_o;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3404_o = n3138_o ? n3334_o : 1'b0;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3406_o = n3138_o ? n3336_o : 1'b0;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3408_o = n3138_o ? n3338_o : 1'b0;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3410_o = n3138_o ? n3340_o : 1'b0;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3412_o = n3138_o ? n3342_o : 1'b0;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3414_o = n3138_o ? n3344_o : 1'b0;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3416_o = n3138_o ? n3347_o : 1'b0;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3418_o = n3138_o ? n3349_o : 1'b0;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3420_o = n3138_o ? n3351_o : 1'b0;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3422_o = n3138_o ? n3353_o : 1'b0;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3424_o = n3138_o ? n3356_o : 1'b0;
  /* control_fsm_rtl.vhd:349:9  */
  assign n3426_o = n3138_o ? n3358_o : 1'b0;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3428_o = n3136_o ? 3'b010 : n3392_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3430_o = n3136_o ? 4'b0000 : n3394_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3432_o = n3136_o ? 3'b001 : n3395_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3434_o = n3136_o ? 4'b0000 : n3397_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3436_o = n3136_o ? 4'b0000 : n3398_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3438_o = n3136_o ? 4'b0000 : n3400_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3441_o = n3136_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3443_o = n3136_o ? 1'b1 : n3402_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3445_o = n3136_o ? 1'b0 : n3404_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3447_o = n3136_o ? 1'b0 : n3406_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3449_o = n3136_o ? 1'b0 : n3408_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3451_o = n3136_o ? 1'b0 : n3410_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3453_o = n3136_o ? 1'b0 : n3412_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3455_o = n3136_o ? 1'b0 : n3414_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3457_o = n3136_o ? 1'b0 : n3416_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3459_o = n3136_o ? 1'b0 : n3418_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3461_o = n3136_o ? 1'b0 : n3420_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3463_o = n3136_o ? 1'b0 : n3422_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3465_o = n3136_o ? 1'b0 : n3424_o;
  /* control_fsm_rtl.vhd:344:9  */
  assign n3467_o = n3136_o ? 1'b0 : n3426_o;
  /* control_fsm_rtl.vhd:444:21  */
  assign n3469_o = state == 3'b001;
  /* control_fsm_rtl.vhd:451:24  */
  assign n3471_o = state == 3'b010;
  /* control_fsm_rtl.vhd:451:13  */
  assign n3474_o = n3471_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:451:13  */
  assign n3477_o = n3471_o ? 3'b101 : 3'b000;
  /* control_fsm_rtl.vhd:451:13  */
  assign n3480_o = n3471_o ? 4'b1101 : 4'b0000;
  /* control_fsm_rtl.vhd:451:13  */
  assign n3483_o = n3471_o ? 4'b1111 : 4'b0000;
  /* control_fsm_rtl.vhd:444:13  */
  assign n3486_o = n3469_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:444:13  */
  assign n3488_o = n3469_o ? 4'b0001 : n3474_o;
  /* control_fsm_rtl.vhd:444:13  */
  assign n3490_o = n3469_o ? 3'b101 : n3477_o;
  /* control_fsm_rtl.vhd:444:13  */
  assign n3492_o = n3469_o ? 4'b1110 : n3480_o;
  /* control_fsm_rtl.vhd:444:13  */
  assign n3494_o = n3469_o ? 4'b1111 : n3483_o;
  /* control_fsm_rtl.vhd:444:13  */
  assign n3497_o = n3469_o ? 2'b10 : 2'b00;
  /* control_fsm_rtl.vhd:443:11  */
  assign n3499_o = s_instr_category == 7'b0000000;
  /* control_fsm_rtl.vhd:462:21  */
  assign n3501_o = state == 3'b001;
  /* control_fsm_rtl.vhd:465:24  */
  assign n3503_o = state == 3'b010;
  /* control_fsm_rtl.vhd:465:13  */
  assign n3506_o = n3503_o ? 6'b100001 : 6'b000000;
  /* control_fsm_rtl.vhd:465:13  */
  assign n3509_o = n3503_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:465:13  */
  assign n3512_o = n3503_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:465:13  */
  assign n3515_o = n3503_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:462:13  */
  assign n3517_o = n3501_o ? 6'b000000 : n3506_o;
  /* control_fsm_rtl.vhd:462:13  */
  assign n3520_o = n3501_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:462:13  */
  assign n3522_o = n3501_o ? 4'b0000 : n3509_o;
  /* control_fsm_rtl.vhd:462:13  */
  assign n3524_o = n3501_o ? 3'b000 : n3512_o;
  /* control_fsm_rtl.vhd:462:13  */
  assign n3526_o = n3501_o ? 4'b0000 : n3515_o;
  /* control_fsm_rtl.vhd:462:13  */
  assign n3529_o = n3501_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:461:11  */
  assign n3531_o = s_instr_category == 7'b0000001;
  /* control_fsm_rtl.vhd:476:21  */
  assign n3533_o = state == 3'b001;
  /* control_fsm_rtl.vhd:479:24  */
  assign n3535_o = state == 3'b010;
  /* control_fsm_rtl.vhd:482:24  */
  assign n3537_o = state == 3'b011;
  /* control_fsm_rtl.vhd:482:13  */
  assign n3540_o = n3537_o ? 6'b100001 : 6'b000000;
  /* control_fsm_rtl.vhd:482:13  */
  assign n3543_o = n3537_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:482:13  */
  assign n3546_o = n3537_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:482:13  */
  assign n3549_o = n3537_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:479:13  */
  assign n3551_o = n3535_o ? 6'b000000 : n3540_o;
  /* control_fsm_rtl.vhd:479:13  */
  assign n3554_o = n3535_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:479:13  */
  assign n3556_o = n3535_o ? 4'b0000 : n3543_o;
  /* control_fsm_rtl.vhd:479:13  */
  assign n3558_o = n3535_o ? 3'b000 : n3546_o;
  /* control_fsm_rtl.vhd:479:13  */
  assign n3560_o = n3535_o ? 4'b0000 : n3549_o;
  /* control_fsm_rtl.vhd:479:13  */
  assign n3563_o = n3535_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:476:13  */
  assign n3565_o = n3533_o ? 6'b000000 : n3551_o;
  /* control_fsm_rtl.vhd:476:13  */
  assign n3567_o = n3533_o ? 3'b010 : n3554_o;
  /* control_fsm_rtl.vhd:476:13  */
  assign n3569_o = n3533_o ? 4'b0001 : n3556_o;
  /* control_fsm_rtl.vhd:476:13  */
  assign n3571_o = n3533_o ? 3'b000 : n3558_o;
  /* control_fsm_rtl.vhd:476:13  */
  assign n3573_o = n3533_o ? 4'b0000 : n3560_o;
  /* control_fsm_rtl.vhd:476:13  */
  assign n3575_o = n3533_o ? 4'b0000 : n3563_o;
  /* control_fsm_rtl.vhd:475:11  */
  assign n3577_o = s_instr_category == 7'b0000010;
  /* control_fsm_rtl.vhd:493:21  */
  assign n3579_o = state == 3'b001;
  /* control_fsm_rtl.vhd:496:24  */
  assign n3581_o = state == 3'b010;
  /* control_fsm_rtl.vhd:496:13  */
  assign n3584_o = n3581_o ? 6'b100001 : 6'b000000;
  /* control_fsm_rtl.vhd:496:13  */
  assign n3587_o = n3581_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:496:13  */
  assign n3590_o = n3581_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:496:13  */
  assign n3593_o = n3581_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:493:13  */
  assign n3595_o = n3579_o ? 6'b000000 : n3584_o;
  /* control_fsm_rtl.vhd:493:13  */
  assign n3598_o = n3579_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:493:13  */
  assign n3600_o = n3579_o ? 4'b0000 : n3587_o;
  /* control_fsm_rtl.vhd:493:13  */
  assign n3602_o = n3579_o ? 3'b000 : n3590_o;
  /* control_fsm_rtl.vhd:493:13  */
  assign n3604_o = n3579_o ? 4'b0000 : n3593_o;
  /* control_fsm_rtl.vhd:493:13  */
  assign n3607_o = n3579_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:492:11  */
  assign n3609_o = s_instr_category == 7'b0000011;
  /* control_fsm_rtl.vhd:507:21  */
  assign n3611_o = state == 3'b001;
  /* control_fsm_rtl.vhd:510:24  */
  assign n3613_o = state == 3'b010;
  /* control_fsm_rtl.vhd:510:13  */
  assign n3616_o = n3613_o ? 6'b100010 : 6'b000000;
  /* control_fsm_rtl.vhd:510:13  */
  assign n3619_o = n3613_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:510:13  */
  assign n3622_o = n3613_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:510:13  */
  assign n3625_o = n3613_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:507:13  */
  assign n3627_o = n3611_o ? 6'b000000 : n3616_o;
  /* control_fsm_rtl.vhd:507:13  */
  assign n3630_o = n3611_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:507:13  */
  assign n3632_o = n3611_o ? 4'b0001 : n3619_o;
  /* control_fsm_rtl.vhd:507:13  */
  assign n3634_o = n3611_o ? 3'b000 : n3622_o;
  /* control_fsm_rtl.vhd:507:13  */
  assign n3636_o = n3611_o ? 4'b0000 : n3625_o;
  /* control_fsm_rtl.vhd:506:11  */
  assign n3638_o = s_instr_category == 7'b0000100;
  /* control_fsm_rtl.vhd:521:21  */
  assign n3640_o = state == 3'b001;
  /* control_fsm_rtl.vhd:524:24  */
  assign n3642_o = state == 3'b010;
  /* control_fsm_rtl.vhd:524:13  */
  assign n3645_o = n3642_o ? 6'b100011 : 6'b000000;
  /* control_fsm_rtl.vhd:524:13  */
  assign n3648_o = n3642_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:524:13  */
  assign n3651_o = n3642_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:524:13  */
  assign n3654_o = n3642_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:521:13  */
  assign n3656_o = n3640_o ? 6'b000000 : n3645_o;
  /* control_fsm_rtl.vhd:521:13  */
  assign n3659_o = n3640_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:521:13  */
  assign n3661_o = n3640_o ? 4'b0000 : n3648_o;
  /* control_fsm_rtl.vhd:521:13  */
  assign n3663_o = n3640_o ? 3'b000 : n3651_o;
  /* control_fsm_rtl.vhd:521:13  */
  assign n3665_o = n3640_o ? 4'b0000 : n3654_o;
  /* control_fsm_rtl.vhd:521:13  */
  assign n3668_o = n3640_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:520:11  */
  assign n3670_o = s_instr_category == 7'b0000101;
  /* control_fsm_rtl.vhd:535:21  */
  assign n3672_o = state == 3'b001;
  /* control_fsm_rtl.vhd:538:24  */
  assign n3674_o = state == 3'b010;
  /* control_fsm_rtl.vhd:541:24  */
  assign n3676_o = state == 3'b011;
  /* control_fsm_rtl.vhd:541:13  */
  assign n3679_o = n3676_o ? 6'b100011 : 6'b000000;
  /* control_fsm_rtl.vhd:541:13  */
  assign n3682_o = n3676_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:541:13  */
  assign n3685_o = n3676_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:541:13  */
  assign n3688_o = n3676_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:538:13  */
  assign n3690_o = n3674_o ? 6'b000000 : n3679_o;
  /* control_fsm_rtl.vhd:538:13  */
  assign n3693_o = n3674_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:538:13  */
  assign n3695_o = n3674_o ? 4'b0000 : n3682_o;
  /* control_fsm_rtl.vhd:538:13  */
  assign n3697_o = n3674_o ? 3'b000 : n3685_o;
  /* control_fsm_rtl.vhd:538:13  */
  assign n3699_o = n3674_o ? 4'b0000 : n3688_o;
  /* control_fsm_rtl.vhd:538:13  */
  assign n3702_o = n3674_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:535:13  */
  assign n3704_o = n3672_o ? 6'b000000 : n3690_o;
  /* control_fsm_rtl.vhd:535:13  */
  assign n3706_o = n3672_o ? 3'b010 : n3693_o;
  /* control_fsm_rtl.vhd:535:13  */
  assign n3708_o = n3672_o ? 4'b0001 : n3695_o;
  /* control_fsm_rtl.vhd:535:13  */
  assign n3710_o = n3672_o ? 3'b000 : n3697_o;
  /* control_fsm_rtl.vhd:535:13  */
  assign n3712_o = n3672_o ? 4'b0000 : n3699_o;
  /* control_fsm_rtl.vhd:535:13  */
  assign n3714_o = n3672_o ? 4'b0000 : n3702_o;
  /* control_fsm_rtl.vhd:534:11  */
  assign n3716_o = s_instr_category == 7'b0000110;
  /* control_fsm_rtl.vhd:552:21  */
  assign n3718_o = state == 3'b001;
  /* control_fsm_rtl.vhd:555:24  */
  assign n3720_o = state == 3'b010;
  /* control_fsm_rtl.vhd:555:13  */
  assign n3723_o = n3720_o ? 6'b100011 : 6'b000000;
  /* control_fsm_rtl.vhd:555:13  */
  assign n3726_o = n3720_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:555:13  */
  assign n3729_o = n3720_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:555:13  */
  assign n3732_o = n3720_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:552:13  */
  assign n3734_o = n3718_o ? 6'b000000 : n3723_o;
  /* control_fsm_rtl.vhd:552:13  */
  assign n3737_o = n3718_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:552:13  */
  assign n3739_o = n3718_o ? 4'b0000 : n3726_o;
  /* control_fsm_rtl.vhd:552:13  */
  assign n3741_o = n3718_o ? 3'b000 : n3729_o;
  /* control_fsm_rtl.vhd:552:13  */
  assign n3743_o = n3718_o ? 4'b0000 : n3732_o;
  /* control_fsm_rtl.vhd:552:13  */
  assign n3746_o = n3718_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:551:11  */
  assign n3748_o = s_instr_category == 7'b0000111;
  /* control_fsm_rtl.vhd:566:21  */
  assign n3750_o = state == 3'b001;
  /* control_fsm_rtl.vhd:569:24  */
  assign n3752_o = state == 3'b010;
  /* control_fsm_rtl.vhd:569:13  */
  assign n3755_o = n3752_o ? 6'b100100 : 6'b000000;
  /* control_fsm_rtl.vhd:569:13  */
  assign n3758_o = n3752_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:569:13  */
  assign n3761_o = n3752_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:569:13  */
  assign n3764_o = n3752_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:566:13  */
  assign n3766_o = n3750_o ? 6'b000000 : n3755_o;
  /* control_fsm_rtl.vhd:566:13  */
  assign n3769_o = n3750_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:566:13  */
  assign n3771_o = n3750_o ? 4'b0001 : n3758_o;
  /* control_fsm_rtl.vhd:566:13  */
  assign n3773_o = n3750_o ? 3'b000 : n3761_o;
  /* control_fsm_rtl.vhd:566:13  */
  assign n3775_o = n3750_o ? 4'b0000 : n3764_o;
  /* control_fsm_rtl.vhd:565:11  */
  assign n3777_o = s_instr_category == 7'b0001000;
  /* control_fsm_rtl.vhd:580:21  */
  assign n3779_o = state == 3'b001;
  /* control_fsm_rtl.vhd:584:24  */
  assign n3781_o = state == 3'b010;
  /* control_fsm_rtl.vhd:584:13  */
  assign n3784_o = n3781_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:580:13  */
  assign n3787_o = n3779_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:580:13  */
  assign n3789_o = n3779_o ? 4'b0001 : n3784_o;
  /* control_fsm_rtl.vhd:580:13  */
  assign n3792_o = n3779_o ? 2'b10 : 2'b00;
  /* control_fsm_rtl.vhd:579:11  */
  assign n3794_o = s_instr_category == 7'b0001001;
  /* control_fsm_rtl.vhd:592:21  */
  assign n3796_o = state == 3'b001;
  /* control_fsm_rtl.vhd:595:24  */
  assign n3798_o = state == 3'b010;
  /* control_fsm_rtl.vhd:595:13  */
  assign n3801_o = n3798_o ? 6'b100101 : 6'b000000;
  /* control_fsm_rtl.vhd:595:13  */
  assign n3804_o = n3798_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:595:13  */
  assign n3807_o = n3798_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:595:13  */
  assign n3810_o = n3798_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:592:13  */
  assign n3812_o = n3796_o ? 6'b000000 : n3801_o;
  /* control_fsm_rtl.vhd:592:13  */
  assign n3815_o = n3796_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:592:13  */
  assign n3817_o = n3796_o ? 4'b0000 : n3804_o;
  /* control_fsm_rtl.vhd:592:13  */
  assign n3819_o = n3796_o ? 3'b000 : n3807_o;
  /* control_fsm_rtl.vhd:592:13  */
  assign n3821_o = n3796_o ? 4'b0000 : n3810_o;
  /* control_fsm_rtl.vhd:592:13  */
  assign n3824_o = n3796_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:591:11  */
  assign n3826_o = s_instr_category == 7'b0001010;
  /* control_fsm_rtl.vhd:606:21  */
  assign n3828_o = state == 3'b001;
  /* control_fsm_rtl.vhd:609:24  */
  assign n3830_o = state == 3'b010;
  /* control_fsm_rtl.vhd:612:24  */
  assign n3832_o = state == 3'b011;
  /* control_fsm_rtl.vhd:612:13  */
  assign n3835_o = n3832_o ? 6'b100101 : 6'b000000;
  /* control_fsm_rtl.vhd:612:13  */
  assign n3838_o = n3832_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:612:13  */
  assign n3841_o = n3832_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:612:13  */
  assign n3844_o = n3832_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:609:13  */
  assign n3846_o = n3830_o ? 6'b000000 : n3835_o;
  /* control_fsm_rtl.vhd:609:13  */
  assign n3849_o = n3830_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:609:13  */
  assign n3851_o = n3830_o ? 4'b0000 : n3838_o;
  /* control_fsm_rtl.vhd:609:13  */
  assign n3853_o = n3830_o ? 3'b000 : n3841_o;
  /* control_fsm_rtl.vhd:609:13  */
  assign n3855_o = n3830_o ? 4'b0000 : n3844_o;
  /* control_fsm_rtl.vhd:609:13  */
  assign n3858_o = n3830_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:606:13  */
  assign n3860_o = n3828_o ? 6'b000000 : n3846_o;
  /* control_fsm_rtl.vhd:606:13  */
  assign n3862_o = n3828_o ? 3'b010 : n3849_o;
  /* control_fsm_rtl.vhd:606:13  */
  assign n3864_o = n3828_o ? 4'b0001 : n3851_o;
  /* control_fsm_rtl.vhd:606:13  */
  assign n3866_o = n3828_o ? 3'b000 : n3853_o;
  /* control_fsm_rtl.vhd:606:13  */
  assign n3868_o = n3828_o ? 4'b0000 : n3855_o;
  /* control_fsm_rtl.vhd:606:13  */
  assign n3870_o = n3828_o ? 4'b0000 : n3858_o;
  /* control_fsm_rtl.vhd:605:11  */
  assign n3872_o = s_instr_category == 7'b0001011;
  /* control_fsm_rtl.vhd:623:21  */
  assign n3874_o = state == 3'b001;
  /* control_fsm_rtl.vhd:626:24  */
  assign n3876_o = state == 3'b010;
  /* control_fsm_rtl.vhd:626:13  */
  assign n3879_o = n3876_o ? 6'b100101 : 6'b000000;
  /* control_fsm_rtl.vhd:626:13  */
  assign n3882_o = n3876_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:626:13  */
  assign n3885_o = n3876_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:626:13  */
  assign n3888_o = n3876_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:623:13  */
  assign n3890_o = n3874_o ? 6'b000000 : n3879_o;
  /* control_fsm_rtl.vhd:623:13  */
  assign n3893_o = n3874_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:623:13  */
  assign n3895_o = n3874_o ? 4'b0000 : n3882_o;
  /* control_fsm_rtl.vhd:623:13  */
  assign n3897_o = n3874_o ? 3'b000 : n3885_o;
  /* control_fsm_rtl.vhd:623:13  */
  assign n3899_o = n3874_o ? 4'b0000 : n3888_o;
  /* control_fsm_rtl.vhd:623:13  */
  assign n3902_o = n3874_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:622:11  */
  assign n3904_o = s_instr_category == 7'b0001100;
  /* control_fsm_rtl.vhd:636:21  */
  assign n3906_o = state == 3'b001;
  /* control_fsm_rtl.vhd:639:24  */
  assign n3908_o = state == 3'b010;
  /* control_fsm_rtl.vhd:639:13  */
  assign n3911_o = n3908_o ? 6'b100110 : 6'b000000;
  /* control_fsm_rtl.vhd:639:13  */
  assign n3914_o = n3908_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:639:13  */
  assign n3917_o = n3908_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:639:13  */
  assign n3920_o = n3908_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:636:13  */
  assign n3922_o = n3906_o ? 6'b000000 : n3911_o;
  /* control_fsm_rtl.vhd:636:13  */
  assign n3925_o = n3906_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:636:13  */
  assign n3927_o = n3906_o ? 4'b0001 : n3914_o;
  /* control_fsm_rtl.vhd:636:13  */
  assign n3929_o = n3906_o ? 3'b000 : n3917_o;
  /* control_fsm_rtl.vhd:636:13  */
  assign n3931_o = n3906_o ? 4'b0000 : n3920_o;
  /* control_fsm_rtl.vhd:635:11  */
  assign n3933_o = s_instr_category == 7'b0001101;
  /* control_fsm_rtl.vhd:650:21  */
  assign n3935_o = state == 3'b001;
  /* control_fsm_rtl.vhd:653:24  */
  assign n3937_o = state == 3'b010;
  /* control_fsm_rtl.vhd:656:24  */
  assign n3939_o = state == 3'b011;
  /* control_fsm_rtl.vhd:656:13  */
  assign n3942_o = n3939_o ? 6'b100101 : 6'b000000;
  /* control_fsm_rtl.vhd:656:13  */
  assign n3945_o = n3939_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:656:13  */
  assign n3948_o = n3939_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:656:13  */
  assign n3951_o = n3939_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:656:13  */
  assign n3954_o = n3939_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:653:13  */
  assign n3956_o = n3937_o ? 6'b000000 : n3942_o;
  /* control_fsm_rtl.vhd:653:13  */
  assign n3959_o = n3937_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:653:13  */
  assign n3961_o = n3937_o ? 4'b0000 : n3945_o;
  /* control_fsm_rtl.vhd:653:13  */
  assign n3963_o = n3937_o ? 3'b000 : n3948_o;
  /* control_fsm_rtl.vhd:653:13  */
  assign n3965_o = n3937_o ? 4'b0000 : n3951_o;
  /* control_fsm_rtl.vhd:653:13  */
  assign n3967_o = n3937_o ? 4'b1000 : n3954_o;
  /* control_fsm_rtl.vhd:650:13  */
  assign n3969_o = n3935_o ? 6'b000000 : n3956_o;
  /* control_fsm_rtl.vhd:650:13  */
  assign n3971_o = n3935_o ? 3'b010 : n3959_o;
  /* control_fsm_rtl.vhd:650:13  */
  assign n3973_o = n3935_o ? 4'b0001 : n3961_o;
  /* control_fsm_rtl.vhd:650:13  */
  assign n3975_o = n3935_o ? 3'b000 : n3963_o;
  /* control_fsm_rtl.vhd:650:13  */
  assign n3977_o = n3935_o ? 4'b0000 : n3965_o;
  /* control_fsm_rtl.vhd:650:13  */
  assign n3979_o = n3935_o ? 4'b0000 : n3967_o;
  /* control_fsm_rtl.vhd:649:11  */
  assign n3981_o = s_instr_category == 7'b0001110;
  /* control_fsm_rtl.vhd:668:21  */
  assign n3983_o = state == 3'b001;
  /* control_fsm_rtl.vhd:671:24  */
  assign n3985_o = state == 3'b010;
  /* control_fsm_rtl.vhd:676:24  */
  assign n3987_o = state == 3'b011;
  /* control_fsm_rtl.vhd:676:13  */
  assign n3990_o = n3987_o ? 6'b100111 : 6'b000000;
  /* control_fsm_rtl.vhd:676:13  */
  assign n3993_o = n3987_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:676:13  */
  assign n3996_o = n3987_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:676:13  */
  assign n3999_o = n3987_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:676:13  */
  assign n4002_o = n3987_o ? 4'b1010 : 4'b0000;
  /* control_fsm_rtl.vhd:671:13  */
  assign n4004_o = n3985_o ? 6'b000000 : n3990_o;
  /* control_fsm_rtl.vhd:671:13  */
  assign n4007_o = n3985_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:671:13  */
  assign n4009_o = n3985_o ? 4'b0001 : n3993_o;
  /* control_fsm_rtl.vhd:671:13  */
  assign n4011_o = n3985_o ? 3'b000 : n3996_o;
  /* control_fsm_rtl.vhd:671:13  */
  assign n4013_o = n3985_o ? 4'b0000 : n3999_o;
  /* control_fsm_rtl.vhd:671:13  */
  assign n4015_o = n3985_o ? 4'b1000 : n4002_o;
  /* control_fsm_rtl.vhd:671:13  */
  assign n4018_o = n3985_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:668:13  */
  assign n4020_o = n3983_o ? 6'b000000 : n4004_o;
  /* control_fsm_rtl.vhd:668:13  */
  assign n4022_o = n3983_o ? 3'b010 : n4007_o;
  /* control_fsm_rtl.vhd:668:13  */
  assign n4024_o = n3983_o ? 4'b0001 : n4009_o;
  /* control_fsm_rtl.vhd:668:13  */
  assign n4026_o = n3983_o ? 3'b000 : n4011_o;
  /* control_fsm_rtl.vhd:668:13  */
  assign n4028_o = n3983_o ? 4'b0000 : n4013_o;
  /* control_fsm_rtl.vhd:668:13  */
  assign n4030_o = n3983_o ? 4'b0000 : n4015_o;
  /* control_fsm_rtl.vhd:668:13  */
  assign n4032_o = n3983_o ? 4'b0000 : n4018_o;
  /* control_fsm_rtl.vhd:667:11  */
  assign n4034_o = s_instr_category == 7'b0001111;
  /* control_fsm_rtl.vhd:688:21  */
  assign n4036_o = state == 3'b001;
  /* control_fsm_rtl.vhd:691:24  */
  assign n4038_o = state == 3'b010;
  /* control_fsm_rtl.vhd:694:24  */
  assign n4040_o = state == 3'b011;
  /* control_fsm_rtl.vhd:694:13  */
  assign n4043_o = n4040_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:694:13  */
  assign n4046_o = n4040_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:694:13  */
  assign n4049_o = n4040_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:691:13  */
  assign n4052_o = n4038_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:691:13  */
  assign n4054_o = n4038_o ? 4'b0000 : n4043_o;
  /* control_fsm_rtl.vhd:691:13  */
  assign n4056_o = n4038_o ? 3'b000 : n4046_o;
  /* control_fsm_rtl.vhd:691:13  */
  assign n4058_o = n4038_o ? 4'b0000 : n4049_o;
  /* control_fsm_rtl.vhd:691:13  */
  assign n4061_o = n4038_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:688:13  */
  assign n4063_o = n4036_o ? 3'b010 : n4052_o;
  /* control_fsm_rtl.vhd:688:13  */
  assign n4065_o = n4036_o ? 4'b0001 : n4054_o;
  /* control_fsm_rtl.vhd:688:13  */
  assign n4067_o = n4036_o ? 3'b000 : n4056_o;
  /* control_fsm_rtl.vhd:688:13  */
  assign n4069_o = n4036_o ? 4'b0000 : n4058_o;
  /* control_fsm_rtl.vhd:688:13  */
  assign n4071_o = n4036_o ? 4'b0000 : n4061_o;
  /* control_fsm_rtl.vhd:687:11  */
  assign n4073_o = s_instr_category == 7'b0010000;
  /* control_fsm_rtl.vhd:704:21  */
  assign n4075_o = state == 3'b001;
  /* control_fsm_rtl.vhd:707:24  */
  assign n4077_o = state == 3'b010;
  /* control_fsm_rtl.vhd:710:24  */
  assign n4079_o = state == 3'b011;
  /* control_fsm_rtl.vhd:710:13  */
  assign n4082_o = n4079_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:710:13  */
  assign n4085_o = n4079_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:710:13  */
  assign n4088_o = n4079_o ? 4'b0010 : 4'b0000;
  /* control_fsm_rtl.vhd:707:13  */
  assign n4091_o = n4077_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:707:13  */
  assign n4093_o = n4077_o ? 4'b0000 : n4082_o;
  /* control_fsm_rtl.vhd:707:13  */
  assign n4095_o = n4077_o ? 3'b000 : n4085_o;
  /* control_fsm_rtl.vhd:707:13  */
  assign n4097_o = n4077_o ? 4'b0000 : n4088_o;
  /* control_fsm_rtl.vhd:707:13  */
  assign n4100_o = n4077_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:704:13  */
  assign n4102_o = n4075_o ? 3'b010 : n4091_o;
  /* control_fsm_rtl.vhd:704:13  */
  assign n4104_o = n4075_o ? 4'b0001 : n4093_o;
  /* control_fsm_rtl.vhd:704:13  */
  assign n4106_o = n4075_o ? 3'b000 : n4095_o;
  /* control_fsm_rtl.vhd:704:13  */
  assign n4108_o = n4075_o ? 4'b0000 : n4097_o;
  /* control_fsm_rtl.vhd:704:13  */
  assign n4110_o = n4075_o ? 4'b0000 : n4100_o;
  /* control_fsm_rtl.vhd:703:11  */
  assign n4112_o = s_instr_category == 7'b0010001;
  /* control_fsm_rtl.vhd:720:21  */
  assign n4114_o = state == 3'b001;
  /* control_fsm_rtl.vhd:723:24  */
  assign n4116_o = state == 3'b010;
  /* control_fsm_rtl.vhd:727:24  */
  assign n4118_o = state == 3'b011;
  /* control_fsm_rtl.vhd:729:38  */
  assign n4119_o = {1'b0, aludata_i};  //  uext
  /* control_fsm_rtl.vhd:729:38  */
  assign n4121_o = n4119_o != 9'b000000000;
  /* control_fsm_rtl.vhd:729:15  */
  assign n4124_o = n4121_o ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:729:15  */
  assign n4127_o = n4121_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:727:13  */
  assign n4130_o = n4118_o ? 6'b111010 : 6'b000000;
  /* control_fsm_rtl.vhd:727:13  */
  assign n4132_o = n4118_o ? n4124_o : 4'b0000;
  /* control_fsm_rtl.vhd:727:13  */
  assign n4135_o = n4118_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:727:13  */
  assign n4137_o = n4118_o ? n4127_o : 4'b0000;
  /* control_fsm_rtl.vhd:727:13  */
  assign n4140_o = n4118_o ? 4'b1011 : 4'b0000;
  /* control_fsm_rtl.vhd:723:13  */
  assign n4142_o = n4116_o ? 6'b000000 : n4130_o;
  /* control_fsm_rtl.vhd:723:13  */
  assign n4145_o = n4116_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:723:13  */
  assign n4147_o = n4116_o ? 4'b0001 : n4132_o;
  /* control_fsm_rtl.vhd:723:13  */
  assign n4149_o = n4116_o ? 3'b000 : n4135_o;
  /* control_fsm_rtl.vhd:723:13  */
  assign n4151_o = n4116_o ? 4'b0000 : n4137_o;
  /* control_fsm_rtl.vhd:723:13  */
  assign n4153_o = n4116_o ? 4'b1000 : n4140_o;
  /* control_fsm_rtl.vhd:720:13  */
  assign n4155_o = n4114_o ? 6'b000000 : n4142_o;
  /* control_fsm_rtl.vhd:720:13  */
  assign n4157_o = n4114_o ? 3'b010 : n4145_o;
  /* control_fsm_rtl.vhd:720:13  */
  assign n4159_o = n4114_o ? 4'b0001 : n4147_o;
  /* control_fsm_rtl.vhd:720:13  */
  assign n4161_o = n4114_o ? 3'b000 : n4149_o;
  /* control_fsm_rtl.vhd:720:13  */
  assign n4163_o = n4114_o ? 4'b0000 : n4151_o;
  /* control_fsm_rtl.vhd:720:13  */
  assign n4165_o = n4114_o ? 4'b0000 : n4153_o;
  /* control_fsm_rtl.vhd:719:11  */
  assign n4167_o = s_instr_category == 7'b0010010;
  /* control_fsm_rtl.vhd:746:21  */
  assign n4169_o = state == 3'b001;
  /* control_fsm_rtl.vhd:749:24  */
  assign n4171_o = state == 3'b010;
  /* control_fsm_rtl.vhd:755:24  */
  assign n4173_o = state == 3'b011;
  /* control_fsm_rtl.vhd:756:25  */
  assign n4174_o = {1'b0, s_help};  //  uext
  /* control_fsm_rtl.vhd:756:25  */
  assign n4176_o = n4174_o != 9'b000000000;
  /* control_fsm_rtl.vhd:756:15  */
  assign n4179_o = n4176_o ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:756:15  */
  assign n4182_o = n4176_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:755:13  */
  assign n4184_o = n4173_o ? n4179_o : 4'b0000;
  /* control_fsm_rtl.vhd:755:13  */
  assign n4187_o = n4173_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:755:13  */
  assign n4189_o = n4173_o ? n4182_o : 4'b0000;
  /* control_fsm_rtl.vhd:755:13  */
  assign n4192_o = n4173_o ? 4'b1011 : 4'b0000;
  /* control_fsm_rtl.vhd:749:13  */
  assign n4195_o = n4171_o ? 6'b111011 : 6'b000000;
  /* control_fsm_rtl.vhd:749:13  */
  assign n4198_o = n4171_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:749:13  */
  assign n4200_o = n4171_o ? 4'b0001 : n4184_o;
  /* control_fsm_rtl.vhd:749:13  */
  assign n4202_o = n4171_o ? 3'b000 : n4187_o;
  /* control_fsm_rtl.vhd:749:13  */
  assign n4204_o = n4171_o ? 4'b0000 : n4189_o;
  /* control_fsm_rtl.vhd:749:13  */
  assign n4206_o = n4171_o ? 4'b0000 : n4192_o;
  /* control_fsm_rtl.vhd:749:13  */
  assign n4209_o = n4171_o ? 4'b0010 : 4'b0000;
  /* control_fsm_rtl.vhd:749:13  */
  assign n4212_o = n4171_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:746:13  */
  assign n4214_o = n4169_o ? 6'b000000 : n4195_o;
  /* control_fsm_rtl.vhd:746:13  */
  assign n4216_o = n4169_o ? 3'b010 : n4198_o;
  /* control_fsm_rtl.vhd:746:13  */
  assign n4218_o = n4169_o ? 4'b0001 : n4200_o;
  /* control_fsm_rtl.vhd:746:13  */
  assign n4220_o = n4169_o ? 3'b000 : n4202_o;
  /* control_fsm_rtl.vhd:746:13  */
  assign n4222_o = n4169_o ? 4'b0000 : n4204_o;
  /* control_fsm_rtl.vhd:746:13  */
  assign n4224_o = n4169_o ? 4'b0000 : n4206_o;
  /* control_fsm_rtl.vhd:746:13  */
  assign n4226_o = n4169_o ? 4'b0000 : n4209_o;
  /* control_fsm_rtl.vhd:746:13  */
  assign n4228_o = n4169_o ? 1'b0 : n4212_o;
  /* control_fsm_rtl.vhd:745:11  */
  assign n4230_o = s_instr_category == 7'b0010011;
  /* control_fsm_rtl.vhd:773:21  */
  assign n4232_o = state == 3'b001;
  /* control_fsm_rtl.vhd:777:24  */
  assign n4234_o = state == 3'b010;
  /* control_fsm_rtl.vhd:783:24  */
  assign n4236_o = state == 3'b011;
  /* control_fsm_rtl.vhd:784:25  */
  assign n4237_o = {1'b0, s_help};  //  uext
  /* control_fsm_rtl.vhd:784:25  */
  assign n4239_o = n4237_o != 9'b000000000;
  /* control_fsm_rtl.vhd:784:15  */
  assign n4242_o = n4239_o ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:784:15  */
  assign n4245_o = n4239_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:783:13  */
  assign n4247_o = n4236_o ? n4242_o : 4'b0000;
  /* control_fsm_rtl.vhd:783:13  */
  assign n4250_o = n4236_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:783:13  */
  assign n4252_o = n4236_o ? n4245_o : 4'b0000;
  /* control_fsm_rtl.vhd:783:13  */
  assign n4255_o = n4236_o ? 4'b1011 : 4'b0000;
  /* control_fsm_rtl.vhd:777:13  */
  assign n4258_o = n4234_o ? 6'b111100 : 6'b000000;
  /* control_fsm_rtl.vhd:777:13  */
  assign n4261_o = n4234_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:777:13  */
  assign n4263_o = n4234_o ? 4'b0001 : n4247_o;
  /* control_fsm_rtl.vhd:777:13  */
  assign n4265_o = n4234_o ? 3'b000 : n4250_o;
  /* control_fsm_rtl.vhd:777:13  */
  assign n4267_o = n4234_o ? 4'b0000 : n4252_o;
  /* control_fsm_rtl.vhd:777:13  */
  assign n4269_o = n4234_o ? 4'b0000 : n4255_o;
  /* control_fsm_rtl.vhd:777:13  */
  assign n4272_o = n4234_o ? 4'b0010 : 4'b0000;
  /* control_fsm_rtl.vhd:777:13  */
  assign n4275_o = n4234_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:773:13  */
  assign n4277_o = n4232_o ? 6'b000000 : n4258_o;
  /* control_fsm_rtl.vhd:773:13  */
  assign n4279_o = n4232_o ? 3'b010 : n4261_o;
  /* control_fsm_rtl.vhd:773:13  */
  assign n4281_o = n4232_o ? 4'b0001 : n4263_o;
  /* control_fsm_rtl.vhd:773:13  */
  assign n4283_o = n4232_o ? 3'b000 : n4265_o;
  /* control_fsm_rtl.vhd:773:13  */
  assign n4285_o = n4232_o ? 4'b0000 : n4267_o;
  /* control_fsm_rtl.vhd:773:13  */
  assign n4287_o = n4232_o ? 4'b0110 : n4269_o;
  /* control_fsm_rtl.vhd:773:13  */
  assign n4289_o = n4232_o ? 4'b0000 : n4272_o;
  /* control_fsm_rtl.vhd:773:13  */
  assign n4291_o = n4232_o ? 1'b0 : n4275_o;
  /* control_fsm_rtl.vhd:772:11  */
  assign n4293_o = s_instr_category == 7'b0010100;
  /* control_fsm_rtl.vhd:801:21  */
  assign n4295_o = state == 3'b001;
  /* control_fsm_rtl.vhd:805:24  */
  assign n4297_o = state == 3'b010;
  /* control_fsm_rtl.vhd:811:24  */
  assign n4299_o = state == 3'b011;
  /* control_fsm_rtl.vhd:812:25  */
  assign n4300_o = {1'b0, s_help};  //  uext
  /* control_fsm_rtl.vhd:812:25  */
  assign n4302_o = n4300_o != 9'b000000000;
  /* control_fsm_rtl.vhd:812:15  */
  assign n4305_o = n4302_o ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:812:15  */
  assign n4308_o = n4302_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:811:13  */
  assign n4310_o = n4299_o ? n4305_o : 4'b0000;
  /* control_fsm_rtl.vhd:811:13  */
  assign n4313_o = n4299_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:811:13  */
  assign n4315_o = n4299_o ? n4308_o : 4'b0000;
  /* control_fsm_rtl.vhd:811:13  */
  assign n4318_o = n4299_o ? 4'b1011 : 4'b0000;
  /* control_fsm_rtl.vhd:805:13  */
  assign n4321_o = n4297_o ? 6'b111100 : 6'b000000;
  /* control_fsm_rtl.vhd:805:13  */
  assign n4324_o = n4297_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:805:13  */
  assign n4326_o = n4297_o ? 4'b0001 : n4310_o;
  /* control_fsm_rtl.vhd:805:13  */
  assign n4328_o = n4297_o ? 3'b000 : n4313_o;
  /* control_fsm_rtl.vhd:805:13  */
  assign n4330_o = n4297_o ? 4'b0000 : n4315_o;
  /* control_fsm_rtl.vhd:805:13  */
  assign n4332_o = n4297_o ? 4'b0000 : n4318_o;
  /* control_fsm_rtl.vhd:805:13  */
  assign n4335_o = n4297_o ? 4'b0010 : 4'b0000;
  /* control_fsm_rtl.vhd:805:13  */
  assign n4338_o = n4297_o ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:801:13  */
  assign n4340_o = n4295_o ? 6'b000000 : n4321_o;
  /* control_fsm_rtl.vhd:801:13  */
  assign n4342_o = n4295_o ? 3'b010 : n4324_o;
  /* control_fsm_rtl.vhd:801:13  */
  assign n4344_o = n4295_o ? 4'b0001 : n4326_o;
  /* control_fsm_rtl.vhd:801:13  */
  assign n4346_o = n4295_o ? 3'b000 : n4328_o;
  /* control_fsm_rtl.vhd:801:13  */
  assign n4348_o = n4295_o ? 4'b0000 : n4330_o;
  /* control_fsm_rtl.vhd:801:13  */
  assign n4350_o = n4295_o ? 4'b0111 : n4332_o;
  /* control_fsm_rtl.vhd:801:13  */
  assign n4352_o = n4295_o ? 4'b0000 : n4335_o;
  /* control_fsm_rtl.vhd:801:13  */
  assign n4354_o = n4295_o ? 1'b0 : n4338_o;
  /* control_fsm_rtl.vhd:800:11  */
  assign n4356_o = s_instr_category == 7'b0010101;
  /* control_fsm_rtl.vhd:828:11  */
  assign n4358_o = s_instr_category == 7'b0010110;
  /* control_fsm_rtl.vhd:836:11  */
  assign n4360_o = s_instr_category == 7'b0010111;
  /* control_fsm_rtl.vhd:846:21  */
  assign n4362_o = state == 3'b001;
  /* control_fsm_rtl.vhd:849:24  */
  assign n4364_o = state == 3'b010;
  /* control_fsm_rtl.vhd:849:13  */
  assign n4367_o = n4364_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:849:13  */
  assign n4370_o = n4364_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:849:13  */
  assign n4373_o = n4364_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:846:13  */
  assign n4376_o = n4362_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:846:13  */
  assign n4378_o = n4362_o ? 4'b0001 : n4367_o;
  /* control_fsm_rtl.vhd:846:13  */
  assign n4380_o = n4362_o ? 3'b000 : n4370_o;
  /* control_fsm_rtl.vhd:846:13  */
  assign n4382_o = n4362_o ? 4'b0000 : n4373_o;
  /* control_fsm_rtl.vhd:845:11  */
  assign n4384_o = s_instr_category == 7'b0011000;
  /* control_fsm_rtl.vhd:859:11  */
  assign n4386_o = s_instr_category == 7'b0011001;
  /* control_fsm_rtl.vhd:868:11  */
  assign n4388_o = s_instr_category == 7'b0011010;
  /* control_fsm_rtl.vhd:878:21  */
  assign n4390_o = state == 3'b001;
  /* control_fsm_rtl.vhd:881:24  */
  assign n4392_o = state == 3'b010;
  /* control_fsm_rtl.vhd:884:24  */
  assign n4394_o = state == 3'b011;
  /* control_fsm_rtl.vhd:884:13  */
  assign n4397_o = n4394_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:884:13  */
  assign n4400_o = n4394_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:884:13  */
  assign n4403_o = n4394_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:884:13  */
  assign n4406_o = n4394_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:881:13  */
  assign n4409_o = n4392_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:881:13  */
  assign n4411_o = n4392_o ? 4'b0000 : n4397_o;
  /* control_fsm_rtl.vhd:881:13  */
  assign n4413_o = n4392_o ? 3'b000 : n4400_o;
  /* control_fsm_rtl.vhd:881:13  */
  assign n4415_o = n4392_o ? 4'b0000 : n4403_o;
  /* control_fsm_rtl.vhd:881:13  */
  assign n4417_o = n4392_o ? 4'b1000 : n4406_o;
  /* control_fsm_rtl.vhd:878:13  */
  assign n4419_o = n4390_o ? 3'b010 : n4409_o;
  /* control_fsm_rtl.vhd:878:13  */
  assign n4421_o = n4390_o ? 4'b0001 : n4411_o;
  /* control_fsm_rtl.vhd:878:13  */
  assign n4423_o = n4390_o ? 3'b000 : n4413_o;
  /* control_fsm_rtl.vhd:878:13  */
  assign n4425_o = n4390_o ? 4'b0000 : n4415_o;
  /* control_fsm_rtl.vhd:878:13  */
  assign n4427_o = n4390_o ? 4'b0000 : n4417_o;
  /* control_fsm_rtl.vhd:877:11  */
  assign n4429_o = s_instr_category == 7'b0011011;
  /* control_fsm_rtl.vhd:896:11  */
  assign n4431_o = s_instr_category == 7'b0011100;
  /* control_fsm_rtl.vhd:905:11  */
  assign n4433_o = s_instr_category == 7'b0011101;
  /* control_fsm_rtl.vhd:915:21  */
  assign n4435_o = state == 3'b001;
  /* control_fsm_rtl.vhd:918:24  */
  assign n4437_o = state == 3'b010;
  /* control_fsm_rtl.vhd:918:13  */
  assign n4440_o = n4437_o ? 6'b111001 : 6'b000000;
  /* control_fsm_rtl.vhd:918:13  */
  assign n4443_o = n4437_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:918:13  */
  assign n4446_o = n4437_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:918:13  */
  assign n4449_o = n4437_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:918:13  */
  assign n4452_o = n4437_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:915:13  */
  assign n4454_o = n4435_o ? 6'b000000 : n4440_o;
  /* control_fsm_rtl.vhd:915:13  */
  assign n4457_o = n4435_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:915:13  */
  assign n4459_o = n4435_o ? 4'b0000 : n4443_o;
  /* control_fsm_rtl.vhd:915:13  */
  assign n4461_o = n4435_o ? 3'b000 : n4446_o;
  /* control_fsm_rtl.vhd:915:13  */
  assign n4463_o = n4435_o ? 4'b0000 : n4449_o;
  /* control_fsm_rtl.vhd:915:13  */
  assign n4465_o = n4435_o ? 4'b0110 : n4452_o;
  /* control_fsm_rtl.vhd:914:11  */
  assign n4467_o = s_instr_category == 7'b0011110;
  /* control_fsm_rtl.vhd:930:21  */
  assign n4469_o = state == 3'b001;
  /* control_fsm_rtl.vhd:933:24  */
  assign n4471_o = state == 3'b010;
  /* control_fsm_rtl.vhd:936:24  */
  assign n4473_o = state == 3'b011;
  /* control_fsm_rtl.vhd:936:13  */
  assign n4476_o = n4473_o ? 6'b111001 : 6'b000000;
  /* control_fsm_rtl.vhd:936:13  */
  assign n4479_o = n4473_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:936:13  */
  assign n4482_o = n4473_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:936:13  */
  assign n4485_o = n4473_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:936:13  */
  assign n4488_o = n4473_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:933:13  */
  assign n4490_o = n4471_o ? 6'b000000 : n4476_o;
  /* control_fsm_rtl.vhd:933:13  */
  assign n4493_o = n4471_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:933:13  */
  assign n4495_o = n4471_o ? 4'b0000 : n4479_o;
  /* control_fsm_rtl.vhd:933:13  */
  assign n4497_o = n4471_o ? 3'b000 : n4482_o;
  /* control_fsm_rtl.vhd:933:13  */
  assign n4499_o = n4471_o ? 4'b0000 : n4485_o;
  /* control_fsm_rtl.vhd:933:13  */
  assign n4501_o = n4471_o ? 4'b1000 : n4488_o;
  /* control_fsm_rtl.vhd:930:13  */
  assign n4503_o = n4469_o ? 6'b000000 : n4490_o;
  /* control_fsm_rtl.vhd:930:13  */
  assign n4505_o = n4469_o ? 3'b010 : n4493_o;
  /* control_fsm_rtl.vhd:930:13  */
  assign n4507_o = n4469_o ? 4'b0001 : n4495_o;
  /* control_fsm_rtl.vhd:930:13  */
  assign n4509_o = n4469_o ? 3'b000 : n4497_o;
  /* control_fsm_rtl.vhd:930:13  */
  assign n4511_o = n4469_o ? 4'b0000 : n4499_o;
  /* control_fsm_rtl.vhd:930:13  */
  assign n4513_o = n4469_o ? 4'b0000 : n4501_o;
  /* control_fsm_rtl.vhd:929:11  */
  assign n4515_o = s_instr_category == 7'b0011111;
  /* control_fsm_rtl.vhd:948:21  */
  assign n4517_o = state == 3'b001;
  /* control_fsm_rtl.vhd:951:24  */
  assign n4519_o = state == 3'b010;
  /* control_fsm_rtl.vhd:951:13  */
  assign n4522_o = n4519_o ? 6'b111001 : 6'b000000;
  /* control_fsm_rtl.vhd:951:13  */
  assign n4525_o = n4519_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:951:13  */
  assign n4528_o = n4519_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:951:13  */
  assign n4531_o = n4519_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:951:13  */
  assign n4534_o = n4519_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:948:13  */
  assign n4536_o = n4517_o ? 6'b000000 : n4522_o;
  /* control_fsm_rtl.vhd:948:13  */
  assign n4539_o = n4517_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:948:13  */
  assign n4541_o = n4517_o ? 4'b0000 : n4525_o;
  /* control_fsm_rtl.vhd:948:13  */
  assign n4543_o = n4517_o ? 3'b000 : n4528_o;
  /* control_fsm_rtl.vhd:948:13  */
  assign n4545_o = n4517_o ? 4'b0000 : n4531_o;
  /* control_fsm_rtl.vhd:948:13  */
  assign n4547_o = n4517_o ? 4'b0111 : n4534_o;
  /* control_fsm_rtl.vhd:947:11  */
  assign n4549_o = s_instr_category == 7'b0100000;
  /* control_fsm_rtl.vhd:963:21  */
  assign n4551_o = state == 3'b001;
  /* control_fsm_rtl.vhd:967:24  */
  assign n4553_o = state == 3'b010;
  /* control_fsm_rtl.vhd:972:24  */
  assign n4555_o = state == 3'b011;
  /* control_fsm_rtl.vhd:972:13  */
  assign n4558_o = n4555_o ? 6'b101011 : 6'b000000;
  /* control_fsm_rtl.vhd:972:13  */
  assign n4561_o = n4555_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:972:13  */
  assign n4564_o = n4555_o ? 3'b111 : 3'b000;
  /* control_fsm_rtl.vhd:972:13  */
  assign n4567_o = n4555_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:972:13  */
  assign n4570_o = n4555_o ? 4'b1100 : 4'b0000;
  /* control_fsm_rtl.vhd:967:13  */
  assign n4572_o = n4553_o ? 6'b101011 : n4558_o;
  /* control_fsm_rtl.vhd:967:13  */
  assign n4575_o = n4553_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:967:13  */
  assign n4577_o = n4553_o ? 4'b0000 : n4561_o;
  /* control_fsm_rtl.vhd:967:13  */
  assign n4579_o = n4553_o ? 3'b000 : n4564_o;
  /* control_fsm_rtl.vhd:967:13  */
  assign n4581_o = n4553_o ? 4'b0011 : n4567_o;
  /* control_fsm_rtl.vhd:967:13  */
  assign n4583_o = n4553_o ? 4'b1100 : n4570_o;
  /* control_fsm_rtl.vhd:963:13  */
  assign n4585_o = n4551_o ? 6'b101011 : n4572_o;
  /* control_fsm_rtl.vhd:963:13  */
  assign n4587_o = n4551_o ? 3'b010 : n4575_o;
  /* control_fsm_rtl.vhd:963:13  */
  assign n4589_o = n4551_o ? 4'b0000 : n4577_o;
  /* control_fsm_rtl.vhd:963:13  */
  assign n4591_o = n4551_o ? 3'b000 : n4579_o;
  /* control_fsm_rtl.vhd:963:13  */
  assign n4593_o = n4551_o ? 4'b0000 : n4581_o;
  /* control_fsm_rtl.vhd:963:13  */
  assign n4595_o = n4551_o ? 4'b1100 : n4583_o;
  /* control_fsm_rtl.vhd:962:11  */
  assign n4597_o = s_instr_category == 7'b0100001;
  /* control_fsm_rtl.vhd:984:21  */
  assign n4599_o = state == 3'b001;
  /* control_fsm_rtl.vhd:989:24  */
  assign n4601_o = state == 3'b010;
  /* control_fsm_rtl.vhd:991:38  */
  assign n4602_o = {1'b0, aludata_i};  //  uext
  /* control_fsm_rtl.vhd:991:38  */
  assign n4604_o = n4602_o != 9'b000000000;
  /* control_fsm_rtl.vhd:991:15  */
  assign n4607_o = n4604_o ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:989:13  */
  assign n4610_o = n4601_o ? 6'b111001 : 6'b000000;
  /* control_fsm_rtl.vhd:989:13  */
  assign n4612_o = n4601_o ? n4607_o : 4'b0000;
  /* control_fsm_rtl.vhd:989:13  */
  assign n4615_o = n4601_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:989:13  */
  assign n4618_o = n4601_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:989:13  */
  assign n4621_o = n4601_o ? 4'b1010 : 4'b0000;
  /* control_fsm_rtl.vhd:984:13  */
  assign n4623_o = n4599_o ? 6'b000000 : n4610_o;
  /* control_fsm_rtl.vhd:984:13  */
  assign n4626_o = n4599_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:984:13  */
  assign n4628_o = n4599_o ? 4'b0001 : n4612_o;
  /* control_fsm_rtl.vhd:984:13  */
  assign n4630_o = n4599_o ? 3'b000 : n4615_o;
  /* control_fsm_rtl.vhd:984:13  */
  assign n4632_o = n4599_o ? 4'b0000 : n4618_o;
  /* control_fsm_rtl.vhd:984:13  */
  assign n4634_o = n4599_o ? 4'b0110 : n4621_o;
  /* control_fsm_rtl.vhd:984:13  */
  assign n4637_o = n4599_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:983:11  */
  assign n4639_o = s_instr_category == 7'b0100010;
  /* control_fsm_rtl.vhd:1008:21  */
  assign n4641_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1011:24  */
  assign n4643_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1016:24  */
  assign n4645_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1018:38  */
  assign n4646_o = {1'b0, aludata_i};  //  uext
  /* control_fsm_rtl.vhd:1018:38  */
  assign n4648_o = n4646_o != 9'b000000000;
  /* control_fsm_rtl.vhd:1018:15  */
  assign n4651_o = n4648_o ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:1016:13  */
  assign n4654_o = n4645_o ? 6'b111001 : 6'b000000;
  /* control_fsm_rtl.vhd:1016:13  */
  assign n4656_o = n4645_o ? n4651_o : 4'b0000;
  /* control_fsm_rtl.vhd:1016:13  */
  assign n4659_o = n4645_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1016:13  */
  assign n4662_o = n4645_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1016:13  */
  assign n4665_o = n4645_o ? 4'b1010 : 4'b0000;
  /* control_fsm_rtl.vhd:1011:13  */
  assign n4667_o = n4643_o ? 6'b000000 : n4654_o;
  /* control_fsm_rtl.vhd:1011:13  */
  assign n4670_o = n4643_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1011:13  */
  assign n4672_o = n4643_o ? 4'b0001 : n4656_o;
  /* control_fsm_rtl.vhd:1011:13  */
  assign n4674_o = n4643_o ? 3'b000 : n4659_o;
  /* control_fsm_rtl.vhd:1011:13  */
  assign n4676_o = n4643_o ? 4'b0000 : n4662_o;
  /* control_fsm_rtl.vhd:1011:13  */
  assign n4678_o = n4643_o ? 4'b1000 : n4665_o;
  /* control_fsm_rtl.vhd:1011:13  */
  assign n4681_o = n4643_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1008:13  */
  assign n4683_o = n4641_o ? 6'b000000 : n4667_o;
  /* control_fsm_rtl.vhd:1008:13  */
  assign n4685_o = n4641_o ? 3'b010 : n4670_o;
  /* control_fsm_rtl.vhd:1008:13  */
  assign n4687_o = n4641_o ? 4'b0001 : n4672_o;
  /* control_fsm_rtl.vhd:1008:13  */
  assign n4689_o = n4641_o ? 3'b000 : n4674_o;
  /* control_fsm_rtl.vhd:1008:13  */
  assign n4691_o = n4641_o ? 4'b0000 : n4676_o;
  /* control_fsm_rtl.vhd:1008:13  */
  assign n4693_o = n4641_o ? 4'b0000 : n4678_o;
  /* control_fsm_rtl.vhd:1008:13  */
  assign n4695_o = n4641_o ? 4'b0000 : n4681_o;
  /* control_fsm_rtl.vhd:1007:11  */
  assign n4697_o = s_instr_category == 7'b0100011;
  /* control_fsm_rtl.vhd:1034:11  */
  assign n4699_o = s_instr_category == 7'b0100100;
  /* control_fsm_rtl.vhd:1044:21  */
  assign n4701_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1047:24  */
  assign n4703_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1047:13  */
  assign n4706_o = n4703_o ? 6'b111111 : 6'b000000;
  /* control_fsm_rtl.vhd:1047:13  */
  assign n4709_o = n4703_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1047:13  */
  assign n4712_o = n4703_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1047:13  */
  assign n4715_o = n4703_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1047:13  */
  assign n4718_o = n4703_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:1044:13  */
  assign n4720_o = n4701_o ? 6'b000000 : n4706_o;
  /* control_fsm_rtl.vhd:1044:13  */
  assign n4723_o = n4701_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1044:13  */
  assign n4725_o = n4701_o ? 4'b0000 : n4709_o;
  /* control_fsm_rtl.vhd:1044:13  */
  assign n4727_o = n4701_o ? 3'b000 : n4712_o;
  /* control_fsm_rtl.vhd:1044:13  */
  assign n4729_o = n4701_o ? 4'b0000 : n4715_o;
  /* control_fsm_rtl.vhd:1044:13  */
  assign n4731_o = n4701_o ? 4'b0110 : n4718_o;
  /* control_fsm_rtl.vhd:1043:11  */
  assign n4733_o = s_instr_category == 7'b0100101;
  /* control_fsm_rtl.vhd:1059:21  */
  assign n4735_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1062:24  */
  assign n4737_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1065:24  */
  assign n4739_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1065:13  */
  assign n4742_o = n4739_o ? 6'b111111 : 6'b000000;
  /* control_fsm_rtl.vhd:1065:13  */
  assign n4745_o = n4739_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1065:13  */
  assign n4748_o = n4739_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1065:13  */
  assign n4751_o = n4739_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1065:13  */
  assign n4754_o = n4739_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1062:13  */
  assign n4756_o = n4737_o ? 6'b000000 : n4742_o;
  /* control_fsm_rtl.vhd:1062:13  */
  assign n4759_o = n4737_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1062:13  */
  assign n4761_o = n4737_o ? 4'b0000 : n4745_o;
  /* control_fsm_rtl.vhd:1062:13  */
  assign n4763_o = n4737_o ? 3'b000 : n4748_o;
  /* control_fsm_rtl.vhd:1062:13  */
  assign n4765_o = n4737_o ? 4'b0000 : n4751_o;
  /* control_fsm_rtl.vhd:1062:13  */
  assign n4767_o = n4737_o ? 4'b1000 : n4754_o;
  /* control_fsm_rtl.vhd:1059:13  */
  assign n4769_o = n4735_o ? 6'b000000 : n4756_o;
  /* control_fsm_rtl.vhd:1059:13  */
  assign n4771_o = n4735_o ? 3'b010 : n4759_o;
  /* control_fsm_rtl.vhd:1059:13  */
  assign n4773_o = n4735_o ? 4'b0001 : n4761_o;
  /* control_fsm_rtl.vhd:1059:13  */
  assign n4775_o = n4735_o ? 3'b000 : n4763_o;
  /* control_fsm_rtl.vhd:1059:13  */
  assign n4777_o = n4735_o ? 4'b0000 : n4765_o;
  /* control_fsm_rtl.vhd:1059:13  */
  assign n4779_o = n4735_o ? 4'b0000 : n4767_o;
  /* control_fsm_rtl.vhd:1058:11  */
  assign n4781_o = s_instr_category == 7'b0100110;
  /* control_fsm_rtl.vhd:1077:21  */
  assign n4783_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1080:24  */
  assign n4785_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1080:13  */
  assign n4788_o = n4785_o ? 6'b111111 : 6'b000000;
  /* control_fsm_rtl.vhd:1080:13  */
  assign n4791_o = n4785_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1080:13  */
  assign n4794_o = n4785_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1080:13  */
  assign n4797_o = n4785_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1080:13  */
  assign n4800_o = n4785_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:1077:13  */
  assign n4802_o = n4783_o ? 6'b000000 : n4788_o;
  /* control_fsm_rtl.vhd:1077:13  */
  assign n4805_o = n4783_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1077:13  */
  assign n4807_o = n4783_o ? 4'b0000 : n4791_o;
  /* control_fsm_rtl.vhd:1077:13  */
  assign n4809_o = n4783_o ? 3'b000 : n4794_o;
  /* control_fsm_rtl.vhd:1077:13  */
  assign n4811_o = n4783_o ? 4'b0000 : n4797_o;
  /* control_fsm_rtl.vhd:1077:13  */
  assign n4813_o = n4783_o ? 4'b0111 : n4800_o;
  /* control_fsm_rtl.vhd:1076:11  */
  assign n4815_o = s_instr_category == 7'b0100111;
  /* control_fsm_rtl.vhd:1092:21  */
  assign n4817_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1095:24  */
  assign n4819_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1102:24  */
  assign n4821_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1105:24  */
  assign n4823_o = state == 3'b100;
  /* control_fsm_rtl.vhd:1106:24  */
  assign n4825_o = s_help == 8'b00000000;
  /* control_fsm_rtl.vhd:1106:15  */
  assign n4828_o = n4825_o ? 6'b111111 : 6'b000000;
  /* control_fsm_rtl.vhd:1106:15  */
  assign n4831_o = n4825_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1106:15  */
  assign n4834_o = n4825_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1106:15  */
  assign n4837_o = n4825_o ? 4'b1110 : 4'b0000;
  /* control_fsm_rtl.vhd:1105:13  */
  assign n4839_o = n4823_o ? n4828_o : 6'b000000;
  /* control_fsm_rtl.vhd:1105:13  */
  assign n4842_o = n4823_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1105:13  */
  assign n4844_o = n4823_o ? n4831_o : 3'b000;
  /* control_fsm_rtl.vhd:1105:13  */
  assign n4846_o = n4823_o ? n4834_o : 4'b0000;
  /* control_fsm_rtl.vhd:1105:13  */
  assign n4848_o = n4823_o ? n4837_o : 4'b0000;
  /* control_fsm_rtl.vhd:1102:13  */
  assign n4850_o = n4821_o ? 6'b000000 : n4839_o;
  /* control_fsm_rtl.vhd:1102:13  */
  assign n4853_o = n4821_o ? 3'b100 : 3'b001;
  /* control_fsm_rtl.vhd:1102:13  */
  assign n4855_o = n4821_o ? 4'b0000 : n4842_o;
  /* control_fsm_rtl.vhd:1102:13  */
  assign n4857_o = n4821_o ? 3'b000 : n4844_o;
  /* control_fsm_rtl.vhd:1102:13  */
  assign n4859_o = n4821_o ? 4'b0000 : n4846_o;
  /* control_fsm_rtl.vhd:1102:13  */
  assign n4861_o = n4821_o ? 4'b1110 : n4848_o;
  /* control_fsm_rtl.vhd:1095:13  */
  assign n4863_o = n4819_o ? 6'b111111 : n4850_o;
  /* control_fsm_rtl.vhd:1095:13  */
  assign n4865_o = n4819_o ? 3'b011 : n4853_o;
  /* control_fsm_rtl.vhd:1095:13  */
  assign n4867_o = n4819_o ? 4'b0000 : n4855_o;
  /* control_fsm_rtl.vhd:1095:13  */
  assign n4869_o = n4819_o ? 3'b100 : n4857_o;
  /* control_fsm_rtl.vhd:1095:13  */
  assign n4871_o = n4819_o ? 4'b0011 : n4859_o;
  /* control_fsm_rtl.vhd:1095:13  */
  assign n4873_o = n4819_o ? 4'b1101 : n4861_o;
  /* control_fsm_rtl.vhd:1095:13  */
  assign n4876_o = n4819_o ? 4'b0010 : 4'b0000;
  /* control_fsm_rtl.vhd:1092:13  */
  assign n4878_o = n4817_o ? 6'b000000 : n4863_o;
  /* control_fsm_rtl.vhd:1092:13  */
  assign n4880_o = n4817_o ? 3'b010 : n4865_o;
  /* control_fsm_rtl.vhd:1092:13  */
  assign n4882_o = n4817_o ? 4'b0000 : n4867_o;
  /* control_fsm_rtl.vhd:1092:13  */
  assign n4884_o = n4817_o ? 3'b000 : n4869_o;
  /* control_fsm_rtl.vhd:1092:13  */
  assign n4886_o = n4817_o ? 4'b0000 : n4871_o;
  /* control_fsm_rtl.vhd:1092:13  */
  assign n4888_o = n4817_o ? 4'b1101 : n4873_o;
  /* control_fsm_rtl.vhd:1092:13  */
  assign n4890_o = n4817_o ? 4'b0000 : n4876_o;
  /* control_fsm_rtl.vhd:1091:11  */
  assign n4892_o = s_instr_category == 7'b0101000;
  /* control_fsm_rtl.vhd:1120:21  */
  assign n4894_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1123:24  */
  assign n4896_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1127:24  */
  assign n4898_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1128:15  */
  assign n4901_o = s_bit_data ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:1127:13  */
  assign n4903_o = n4898_o ? n4901_o : 4'b0000;
  /* control_fsm_rtl.vhd:1123:13  */
  assign n4906_o = n4896_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1123:13  */
  assign n4908_o = n4896_o ? 4'b0001 : n4903_o;
  /* control_fsm_rtl.vhd:1123:13  */
  assign n4911_o = n4896_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1120:13  */
  assign n4913_o = n4894_o ? 3'b010 : n4906_o;
  /* control_fsm_rtl.vhd:1120:13  */
  assign n4915_o = n4894_o ? 4'b0001 : n4908_o;
  /* control_fsm_rtl.vhd:1120:13  */
  assign n4917_o = n4894_o ? 4'b0000 : n4911_o;
  /* control_fsm_rtl.vhd:1119:11  */
  assign n4919_o = s_instr_category == 7'b0101001;
  /* control_fsm_rtl.vhd:1139:21  */
  assign n4921_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1142:24  */
  assign n4923_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1147:24  */
  assign n4925_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1151:15  */
  assign n4928_o = s_bit_data ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:1147:13  */
  assign n4930_o = n4925_o ? n4928_o : 4'b0000;
  /* control_fsm_rtl.vhd:1147:13  */
  assign n4933_o = n4925_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:1147:13  */
  assign n4936_o = n4925_o ? 4'b1010 : 4'b0000;
  /* control_fsm_rtl.vhd:1142:13  */
  assign n4939_o = n4923_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1142:13  */
  assign n4941_o = n4923_o ? 4'b0001 : n4930_o;
  /* control_fsm_rtl.vhd:1142:13  */
  assign n4943_o = n4923_o ? 3'b000 : n4933_o;
  /* control_fsm_rtl.vhd:1142:13  */
  assign n4945_o = n4923_o ? 4'b1000 : n4936_o;
  /* control_fsm_rtl.vhd:1142:13  */
  assign n4948_o = n4923_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1139:13  */
  assign n4950_o = n4921_o ? 3'b010 : n4939_o;
  /* control_fsm_rtl.vhd:1139:13  */
  assign n4952_o = n4921_o ? 4'b0001 : n4941_o;
  /* control_fsm_rtl.vhd:1139:13  */
  assign n4954_o = n4921_o ? 3'b000 : n4943_o;
  /* control_fsm_rtl.vhd:1139:13  */
  assign n4956_o = n4921_o ? 4'b0000 : n4945_o;
  /* control_fsm_rtl.vhd:1139:13  */
  assign n4958_o = n4921_o ? 4'b0000 : n4948_o;
  /* control_fsm_rtl.vhd:1138:11  */
  assign n4960_o = s_instr_category == 7'b0101010;
  /* control_fsm_rtl.vhd:1162:21  */
  assign n4962_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1165:24  */
  assign n4964_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1166:15  */
  assign n4967_o = n2628_o ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:1165:13  */
  assign n4969_o = n4964_o ? n4967_o : 4'b0000;
  /* control_fsm_rtl.vhd:1162:13  */
  assign n4972_o = n4962_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1162:13  */
  assign n4974_o = n4962_o ? 4'b0001 : n4969_o;
  /* control_fsm_rtl.vhd:1161:11  */
  assign n4976_o = s_instr_category == 7'b0101011;
  /* control_fsm_rtl.vhd:1176:11  */
  assign n4978_o = s_instr_category == 7'b0101100;
  /* control_fsm_rtl.vhd:1183:21  */
  assign n4980_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1186:24  */
  assign n4982_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1190:24  */
  assign n4984_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1191:29  */
  assign n4985_o = ~s_bit_data;
  /* control_fsm_rtl.vhd:1191:15  */
  assign n4988_o = n4985_o ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:1190:13  */
  assign n4990_o = n4984_o ? n4988_o : 4'b0000;
  /* control_fsm_rtl.vhd:1186:13  */
  assign n4993_o = n4982_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1186:13  */
  assign n4995_o = n4982_o ? 4'b0001 : n4990_o;
  /* control_fsm_rtl.vhd:1186:13  */
  assign n4998_o = n4982_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1183:13  */
  assign n5000_o = n4980_o ? 3'b010 : n4993_o;
  /* control_fsm_rtl.vhd:1183:13  */
  assign n5002_o = n4980_o ? 4'b0001 : n4995_o;
  /* control_fsm_rtl.vhd:1183:13  */
  assign n5004_o = n4980_o ? 4'b0000 : n4998_o;
  /* control_fsm_rtl.vhd:1182:11  */
  assign n5006_o = s_instr_category == 7'b0101101;
  /* control_fsm_rtl.vhd:1202:21  */
  assign n5008_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1205:24  */
  assign n5010_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1206:21  */
  assign n5011_o = ~n2628_o;
  /* control_fsm_rtl.vhd:1206:15  */
  assign n5014_o = n5011_o ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:1205:13  */
  assign n5016_o = n5010_o ? n5014_o : 4'b0000;
  /* control_fsm_rtl.vhd:1202:13  */
  assign n5019_o = n5008_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1202:13  */
  assign n5021_o = n5008_o ? 4'b0001 : n5016_o;
  /* control_fsm_rtl.vhd:1201:11  */
  assign n5023_o = s_instr_category == 7'b0101110;
  /* control_fsm_rtl.vhd:1217:21  */
  assign n5025_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1220:24  */
  assign n5027_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1221:32  */
  assign n5029_o = acc != 8'b00000000;
  /* control_fsm_rtl.vhd:1221:15  */
  assign n5032_o = n5029_o ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:1220:13  */
  assign n5034_o = n5027_o ? n5032_o : 4'b0000;
  /* control_fsm_rtl.vhd:1217:13  */
  assign n5037_o = n5025_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1217:13  */
  assign n5039_o = n5025_o ? 4'b0001 : n5034_o;
  /* control_fsm_rtl.vhd:1216:11  */
  assign n5041_o = s_instr_category == 7'b0101111;
  /* control_fsm_rtl.vhd:1232:21  */
  assign n5043_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1235:24  */
  assign n5045_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1236:32  */
  assign n5047_o = acc == 8'b00000000;
  /* control_fsm_rtl.vhd:1236:15  */
  assign n5050_o = n5047_o ? 4'b0010 : 4'b0001;
  /* control_fsm_rtl.vhd:1235:13  */
  assign n5052_o = n5045_o ? n5050_o : 4'b0000;
  /* control_fsm_rtl.vhd:1232:13  */
  assign n5055_o = n5043_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1232:13  */
  assign n5057_o = n5043_o ? 4'b0001 : n5052_o;
  /* control_fsm_rtl.vhd:1231:11  */
  assign n5059_o = s_instr_category == 7'b0110000;
  /* control_fsm_rtl.vhd:1247:21  */
  assign n5061_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1252:24  */
  assign n5063_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1259:24  */
  assign n5065_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1259:13  */
  assign n5068_o = n5065_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:1259:13  */
  assign n5071_o = n5065_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1259:13  */
  assign n5074_o = n5065_o ? 4'b1101 : 4'b0000;
  /* control_fsm_rtl.vhd:1259:13  */
  assign n5077_o = n5065_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:1252:13  */
  assign n5080_o = n5063_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1252:13  */
  assign n5082_o = n5063_o ? 4'b0001 : n5068_o;
  /* control_fsm_rtl.vhd:1252:13  */
  assign n5084_o = n5063_o ? 3'b101 : n5071_o;
  /* control_fsm_rtl.vhd:1252:13  */
  assign n5086_o = n5063_o ? 4'b1100 : n5074_o;
  /* control_fsm_rtl.vhd:1252:13  */
  assign n5088_o = n5063_o ? 4'b0101 : n5077_o;
  /* control_fsm_rtl.vhd:1252:13  */
  assign n5091_o = n5063_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1247:13  */
  assign n5093_o = n5061_o ? 3'b010 : n5080_o;
  /* control_fsm_rtl.vhd:1247:13  */
  assign n5095_o = n5061_o ? 4'b0001 : n5082_o;
  /* control_fsm_rtl.vhd:1247:13  */
  assign n5097_o = n5061_o ? 3'b001 : n5084_o;
  /* control_fsm_rtl.vhd:1247:13  */
  assign n5099_o = n5061_o ? 4'b0000 : n5086_o;
  /* control_fsm_rtl.vhd:1247:13  */
  assign n5101_o = n5061_o ? 4'b0000 : n5088_o;
  /* control_fsm_rtl.vhd:1247:13  */
  assign n5103_o = n5061_o ? 4'b0000 : n5091_o;
  /* control_fsm_rtl.vhd:1247:13  */
  assign n5106_o = n5061_o ? 2'b01 : 2'b00;
  /* control_fsm_rtl.vhd:1246:11  */
  assign n5108_o = s_instr_category == 7'b0110001;
  /* control_fsm_rtl.vhd:1270:21  */
  assign n5110_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1273:24  */
  assign n5112_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1277:24  */
  assign n5114_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1277:13  */
  assign n5117_o = n5114_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:1273:13  */
  assign n5120_o = n5112_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1273:13  */
  assign n5122_o = n5112_o ? 4'b0001 : n5117_o;
  /* control_fsm_rtl.vhd:1273:13  */
  assign n5125_o = n5112_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1270:13  */
  assign n5127_o = n5110_o ? 3'b010 : n5120_o;
  /* control_fsm_rtl.vhd:1270:13  */
  assign n5129_o = n5110_o ? 4'b0001 : n5122_o;
  /* control_fsm_rtl.vhd:1270:13  */
  assign n5131_o = n5110_o ? 4'b0000 : n5125_o;
  /* control_fsm_rtl.vhd:1269:11  */
  assign n5133_o = s_instr_category == 7'b0110010;
  /* control_fsm_rtl.vhd:1285:21  */
  assign n5135_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1288:24  */
  assign n5137_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1288:13  */
  assign n5140_o = n5137_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1288:13  */
  assign n5143_o = n5137_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1288:13  */
  assign n5146_o = n5137_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1285:13  */
  assign n5149_o = n5135_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1285:13  */
  assign n5151_o = n5135_o ? 4'b0000 : n5140_o;
  /* control_fsm_rtl.vhd:1285:13  */
  assign n5153_o = n5135_o ? 3'b000 : n5143_o;
  /* control_fsm_rtl.vhd:1285:13  */
  assign n5155_o = n5135_o ? 4'b0000 : n5146_o;
  /* control_fsm_rtl.vhd:1285:13  */
  assign n5158_o = n5135_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:1284:11  */
  assign n5160_o = s_instr_category == 7'b0110011;
  /* control_fsm_rtl.vhd:1297:21  */
  assign n5162_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1300:24  */
  assign n5164_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1303:24  */
  assign n5166_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1303:13  */
  assign n5169_o = n5166_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1303:13  */
  assign n5172_o = n5166_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1303:13  */
  assign n5175_o = n5166_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1300:13  */
  assign n5178_o = n5164_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1300:13  */
  assign n5180_o = n5164_o ? 4'b0000 : n5169_o;
  /* control_fsm_rtl.vhd:1300:13  */
  assign n5182_o = n5164_o ? 3'b000 : n5172_o;
  /* control_fsm_rtl.vhd:1300:13  */
  assign n5184_o = n5164_o ? 4'b0000 : n5175_o;
  /* control_fsm_rtl.vhd:1300:13  */
  assign n5187_o = n5164_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1297:13  */
  assign n5189_o = n5162_o ? 3'b010 : n5178_o;
  /* control_fsm_rtl.vhd:1297:13  */
  assign n5191_o = n5162_o ? 4'b0001 : n5180_o;
  /* control_fsm_rtl.vhd:1297:13  */
  assign n5193_o = n5162_o ? 3'b000 : n5182_o;
  /* control_fsm_rtl.vhd:1297:13  */
  assign n5195_o = n5162_o ? 4'b0000 : n5184_o;
  /* control_fsm_rtl.vhd:1297:13  */
  assign n5197_o = n5162_o ? 4'b0000 : n5187_o;
  /* control_fsm_rtl.vhd:1296:11  */
  assign n5199_o = s_instr_category == 7'b0110100;
  /* control_fsm_rtl.vhd:1313:21  */
  assign n5201_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1316:24  */
  assign n5203_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1316:13  */
  assign n5206_o = n5203_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1316:13  */
  assign n5209_o = n5203_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1316:13  */
  assign n5212_o = n5203_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1313:13  */
  assign n5215_o = n5201_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1313:13  */
  assign n5217_o = n5201_o ? 4'b0000 : n5206_o;
  /* control_fsm_rtl.vhd:1313:13  */
  assign n5219_o = n5201_o ? 3'b000 : n5209_o;
  /* control_fsm_rtl.vhd:1313:13  */
  assign n5221_o = n5201_o ? 4'b0000 : n5212_o;
  /* control_fsm_rtl.vhd:1313:13  */
  assign n5224_o = n5201_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:1312:11  */
  assign n5226_o = s_instr_category == 7'b0110101;
  /* control_fsm_rtl.vhd:1326:21  */
  assign n5228_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1329:24  */
  assign n5230_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1329:13  */
  assign n5233_o = n5230_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1329:13  */
  assign n5236_o = n5230_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1329:13  */
  assign n5239_o = n5230_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:1326:13  */
  assign n5242_o = n5228_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1326:13  */
  assign n5244_o = n5228_o ? 4'b0001 : n5233_o;
  /* control_fsm_rtl.vhd:1326:13  */
  assign n5246_o = n5228_o ? 3'b000 : n5236_o;
  /* control_fsm_rtl.vhd:1326:13  */
  assign n5248_o = n5228_o ? 4'b0000 : n5239_o;
  /* control_fsm_rtl.vhd:1325:11  */
  assign n5250_o = s_instr_category == 7'b0110110;
  /* control_fsm_rtl.vhd:1338:11  */
  assign n5252_o = s_instr_category == 7'b0110111;
  /* control_fsm_rtl.vhd:1348:21  */
  assign n5254_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1352:24  */
  assign n5256_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1355:24  */
  assign n5258_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1355:13  */
  assign n5261_o = n5258_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1355:13  */
  assign n5264_o = n5258_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1355:13  */
  assign n5267_o = n5258_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1355:13  */
  assign n5270_o = n5258_o ? 4'b1010 : 4'b0000;
  /* control_fsm_rtl.vhd:1352:13  */
  assign n5273_o = n5256_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1352:13  */
  assign n5275_o = n5256_o ? 4'b0000 : n5261_o;
  /* control_fsm_rtl.vhd:1352:13  */
  assign n5277_o = n5256_o ? 3'b000 : n5264_o;
  /* control_fsm_rtl.vhd:1352:13  */
  assign n5279_o = n5256_o ? 4'b0000 : n5267_o;
  /* control_fsm_rtl.vhd:1352:13  */
  assign n5281_o = n5256_o ? 4'b1000 : n5270_o;
  /* control_fsm_rtl.vhd:1348:13  */
  assign n5283_o = n5254_o ? 3'b010 : n5273_o;
  /* control_fsm_rtl.vhd:1348:13  */
  assign n5285_o = n5254_o ? 4'b0001 : n5275_o;
  /* control_fsm_rtl.vhd:1348:13  */
  assign n5287_o = n5254_o ? 3'b000 : n5277_o;
  /* control_fsm_rtl.vhd:1348:13  */
  assign n5289_o = n5254_o ? 4'b0000 : n5279_o;
  /* control_fsm_rtl.vhd:1348:13  */
  assign n5291_o = n5254_o ? 4'b0000 : n5281_o;
  /* control_fsm_rtl.vhd:1348:13  */
  assign n5294_o = n5254_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1347:11  */
  assign n5296_o = s_instr_category == 7'b0111000;
  /* control_fsm_rtl.vhd:1366:21  */
  assign n5298_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1370:24  */
  assign n5300_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1370:13  */
  assign n5303_o = n5300_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1370:13  */
  assign n5306_o = n5300_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1370:13  */
  assign n5309_o = n5300_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:1370:13  */
  assign n5312_o = n5300_o ? 4'b1010 : 4'b0000;
  /* control_fsm_rtl.vhd:1366:13  */
  assign n5315_o = n5298_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1366:13  */
  assign n5317_o = n5298_o ? 4'b0001 : n5303_o;
  /* control_fsm_rtl.vhd:1366:13  */
  assign n5319_o = n5298_o ? 3'b000 : n5306_o;
  /* control_fsm_rtl.vhd:1366:13  */
  assign n5321_o = n5298_o ? 4'b0000 : n5309_o;
  /* control_fsm_rtl.vhd:1366:13  */
  assign n5323_o = n5298_o ? 4'b0000 : n5312_o;
  /* control_fsm_rtl.vhd:1366:13  */
  assign n5326_o = n5298_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1365:11  */
  assign n5328_o = s_instr_category == 7'b0111001;
  /* control_fsm_rtl.vhd:1381:21  */
  assign n5330_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1384:24  */
  assign n5332_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1384:13  */
  assign n5335_o = n5332_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1384:13  */
  assign n5338_o = n5332_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1384:13  */
  assign n5341_o = n5332_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:1384:13  */
  assign n5344_o = n5332_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1381:13  */
  assign n5347_o = n5330_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1381:13  */
  assign n5349_o = n5330_o ? 4'b0001 : n5335_o;
  /* control_fsm_rtl.vhd:1381:13  */
  assign n5351_o = n5330_o ? 3'b000 : n5338_o;
  /* control_fsm_rtl.vhd:1381:13  */
  assign n5353_o = n5330_o ? 4'b0000 : n5341_o;
  /* control_fsm_rtl.vhd:1381:13  */
  assign n5355_o = n5330_o ? 4'b0000 : n5344_o;
  /* control_fsm_rtl.vhd:1380:11  */
  assign n5357_o = s_instr_category == 7'b0111010;
  /* control_fsm_rtl.vhd:1395:21  */
  assign n5359_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1399:24  */
  assign n5361_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1399:13  */
  assign n5364_o = n5361_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1399:13  */
  assign n5367_o = n5361_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1399:13  */
  assign n5370_o = n5361_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1399:13  */
  assign n5373_o = n5361_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1395:13  */
  assign n5376_o = n5359_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1395:13  */
  assign n5378_o = n5359_o ? 4'b0001 : n5364_o;
  /* control_fsm_rtl.vhd:1395:13  */
  assign n5380_o = n5359_o ? 3'b000 : n5367_o;
  /* control_fsm_rtl.vhd:1395:13  */
  assign n5382_o = n5359_o ? 4'b0000 : n5370_o;
  /* control_fsm_rtl.vhd:1395:13  */
  assign n5384_o = n5359_o ? 4'b0110 : n5373_o;
  /* control_fsm_rtl.vhd:1394:11  */
  assign n5386_o = s_instr_category == 7'b0111011;
  /* control_fsm_rtl.vhd:1410:21  */
  assign n5388_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1413:24  */
  assign n5390_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1417:24  */
  assign n5392_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1417:13  */
  assign n5395_o = n5392_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1417:13  */
  assign n5398_o = n5392_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1417:13  */
  assign n5401_o = n5392_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1417:13  */
  assign n5404_o = n5392_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1413:13  */
  assign n5407_o = n5390_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1413:13  */
  assign n5409_o = n5390_o ? 4'b0001 : n5395_o;
  /* control_fsm_rtl.vhd:1413:13  */
  assign n5411_o = n5390_o ? 3'b000 : n5398_o;
  /* control_fsm_rtl.vhd:1413:13  */
  assign n5413_o = n5390_o ? 4'b0000 : n5401_o;
  /* control_fsm_rtl.vhd:1413:13  */
  assign n5415_o = n5390_o ? 4'b1000 : n5404_o;
  /* control_fsm_rtl.vhd:1410:13  */
  assign n5417_o = n5388_o ? 3'b010 : n5407_o;
  /* control_fsm_rtl.vhd:1410:13  */
  assign n5419_o = n5388_o ? 4'b0001 : n5409_o;
  /* control_fsm_rtl.vhd:1410:13  */
  assign n5421_o = n5388_o ? 3'b000 : n5411_o;
  /* control_fsm_rtl.vhd:1410:13  */
  assign n5423_o = n5388_o ? 4'b0000 : n5413_o;
  /* control_fsm_rtl.vhd:1410:13  */
  assign n5425_o = n5388_o ? 4'b0000 : n5415_o;
  /* control_fsm_rtl.vhd:1409:11  */
  assign n5427_o = s_instr_category == 7'b0111100;
  /* control_fsm_rtl.vhd:1428:21  */
  assign n5429_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1432:24  */
  assign n5431_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1432:13  */
  assign n5434_o = n5431_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1432:13  */
  assign n5437_o = n5431_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1432:13  */
  assign n5440_o = n5431_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1432:13  */
  assign n5443_o = n5431_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1428:13  */
  assign n5446_o = n5429_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1428:13  */
  assign n5448_o = n5429_o ? 4'b0001 : n5434_o;
  /* control_fsm_rtl.vhd:1428:13  */
  assign n5450_o = n5429_o ? 3'b000 : n5437_o;
  /* control_fsm_rtl.vhd:1428:13  */
  assign n5452_o = n5429_o ? 4'b0000 : n5440_o;
  /* control_fsm_rtl.vhd:1428:13  */
  assign n5454_o = n5429_o ? 4'b0111 : n5443_o;
  /* control_fsm_rtl.vhd:1427:11  */
  assign n5456_o = s_instr_category == 7'b0111101;
  /* control_fsm_rtl.vhd:1443:21  */
  assign n5458_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1446:24  */
  assign n5460_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1450:24  */
  assign n5462_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1450:13  */
  assign n5465_o = n5462_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1450:13  */
  assign n5468_o = n5462_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1450:13  */
  assign n5471_o = n5462_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:1450:13  */
  assign n5474_o = n5462_o ? 4'b1010 : 4'b0000;
  /* control_fsm_rtl.vhd:1446:13  */
  assign n5477_o = n5460_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1446:13  */
  assign n5479_o = n5460_o ? 4'b0001 : n5465_o;
  /* control_fsm_rtl.vhd:1446:13  */
  assign n5481_o = n5460_o ? 3'b000 : n5468_o;
  /* control_fsm_rtl.vhd:1446:13  */
  assign n5483_o = n5460_o ? 4'b0000 : n5471_o;
  /* control_fsm_rtl.vhd:1446:13  */
  assign n5485_o = n5460_o ? 4'b0000 : n5474_o;
  /* control_fsm_rtl.vhd:1446:13  */
  assign n5488_o = n5460_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1443:13  */
  assign n5490_o = n5458_o ? 3'b010 : n5477_o;
  /* control_fsm_rtl.vhd:1443:13  */
  assign n5492_o = n5458_o ? 4'b0001 : n5479_o;
  /* control_fsm_rtl.vhd:1443:13  */
  assign n5494_o = n5458_o ? 3'b000 : n5481_o;
  /* control_fsm_rtl.vhd:1443:13  */
  assign n5496_o = n5458_o ? 4'b0000 : n5483_o;
  /* control_fsm_rtl.vhd:1443:13  */
  assign n5498_o = n5458_o ? 4'b0000 : n5485_o;
  /* control_fsm_rtl.vhd:1443:13  */
  assign n5500_o = n5458_o ? 4'b0000 : n5488_o;
  /* control_fsm_rtl.vhd:1442:11  */
  assign n5502_o = s_instr_category == 7'b0111110;
  /* control_fsm_rtl.vhd:1460:11  */
  assign n5504_o = s_instr_category == 7'b0111111;
  /* control_fsm_rtl.vhd:1470:21  */
  assign n5506_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1473:24  */
  assign n5508_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1476:24  */
  assign n5510_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1476:13  */
  assign n5513_o = n5510_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1476:13  */
  assign n5516_o = n5510_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1476:13  */
  assign n5519_o = n5510_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1476:13  */
  assign n5522_o = n5510_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:1473:13  */
  assign n5525_o = n5508_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1473:13  */
  assign n5527_o = n5508_o ? 4'b0000 : n5513_o;
  /* control_fsm_rtl.vhd:1473:13  */
  assign n5529_o = n5508_o ? 3'b000 : n5516_o;
  /* control_fsm_rtl.vhd:1473:13  */
  assign n5531_o = n5508_o ? 4'b0000 : n5519_o;
  /* control_fsm_rtl.vhd:1473:13  */
  assign n5533_o = n5508_o ? 4'b1000 : n5522_o;
  /* control_fsm_rtl.vhd:1470:13  */
  assign n5535_o = n5506_o ? 3'b010 : n5525_o;
  /* control_fsm_rtl.vhd:1470:13  */
  assign n5537_o = n5506_o ? 4'b0001 : n5527_o;
  /* control_fsm_rtl.vhd:1470:13  */
  assign n5539_o = n5506_o ? 3'b000 : n5529_o;
  /* control_fsm_rtl.vhd:1470:13  */
  assign n5541_o = n5506_o ? 4'b0000 : n5531_o;
  /* control_fsm_rtl.vhd:1470:13  */
  assign n5543_o = n5506_o ? 4'b0000 : n5533_o;
  /* control_fsm_rtl.vhd:1469:11  */
  assign n5545_o = s_instr_category == 7'b1000000;
  /* control_fsm_rtl.vhd:1487:21  */
  assign n5547_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1490:24  */
  assign n5549_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1490:13  */
  assign n5552_o = n5549_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1490:13  */
  assign n5555_o = n5549_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1490:13  */
  assign n5558_o = n5549_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:1490:13  */
  assign n5561_o = n5549_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:1487:13  */
  assign n5564_o = n5547_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1487:13  */
  assign n5566_o = n5547_o ? 4'b0001 : n5552_o;
  /* control_fsm_rtl.vhd:1487:13  */
  assign n5568_o = n5547_o ? 3'b000 : n5555_o;
  /* control_fsm_rtl.vhd:1487:13  */
  assign n5570_o = n5547_o ? 4'b0000 : n5558_o;
  /* control_fsm_rtl.vhd:1487:13  */
  assign n5572_o = n5547_o ? 4'b0000 : n5561_o;
  /* control_fsm_rtl.vhd:1486:11  */
  assign n5574_o = s_instr_category == 7'b1000001;
  /* control_fsm_rtl.vhd:1501:21  */
  assign n5576_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1505:24  */
  assign n5578_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1505:13  */
  assign n5581_o = n5578_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:1505:13  */
  assign n5584_o = n5578_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1505:13  */
  assign n5587_o = n5578_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:1501:13  */
  assign n5590_o = n5576_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1501:13  */
  assign n5592_o = n5576_o ? 4'b0101 : n5581_o;
  /* control_fsm_rtl.vhd:1501:13  */
  assign n5594_o = n5576_o ? 3'b000 : n5584_o;
  /* control_fsm_rtl.vhd:1501:13  */
  assign n5596_o = n5576_o ? 4'b0000 : n5587_o;
  /* control_fsm_rtl.vhd:1501:13  */
  assign n5599_o = n5576_o ? 2'b11 : 2'b00;
  /* control_fsm_rtl.vhd:1500:11  */
  assign n5601_o = s_instr_category == 7'b1000010;
  /* control_fsm_rtl.vhd:1515:21  */
  assign n5603_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1519:24  */
  assign n5605_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1519:13  */
  assign n5608_o = n5605_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:1519:13  */
  assign n5611_o = n5605_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1519:13  */
  assign n5614_o = n5605_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:1515:13  */
  assign n5617_o = n5603_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1515:13  */
  assign n5619_o = n5603_o ? 4'b1001 : n5608_o;
  /* control_fsm_rtl.vhd:1515:13  */
  assign n5621_o = n5603_o ? 3'b000 : n5611_o;
  /* control_fsm_rtl.vhd:1515:13  */
  assign n5623_o = n5603_o ? 4'b0000 : n5614_o;
  /* control_fsm_rtl.vhd:1515:13  */
  assign n5626_o = n5603_o ? 2'b11 : 2'b00;
  /* control_fsm_rtl.vhd:1514:11  */
  assign n5628_o = s_instr_category == 7'b1000011;
  /* control_fsm_rtl.vhd:1529:21  */
  assign n5630_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1532:24  */
  assign n5632_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1532:13  */
  assign n5635_o = n5632_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1532:13  */
  assign n5638_o = n5632_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1532:13  */
  assign n5641_o = n5632_o ? 4'b1111 : 4'b0000;
  /* control_fsm_rtl.vhd:1529:13  */
  assign n5644_o = n5630_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1529:13  */
  assign n5646_o = n5630_o ? 4'b0000 : n5635_o;
  /* control_fsm_rtl.vhd:1529:13  */
  assign n5648_o = n5630_o ? 3'b000 : n5638_o;
  /* control_fsm_rtl.vhd:1529:13  */
  assign n5650_o = n5630_o ? 4'b0000 : n5641_o;
  /* control_fsm_rtl.vhd:1529:13  */
  assign n5653_o = n5630_o ? 2'b10 : 2'b00;
  /* control_fsm_rtl.vhd:1528:11  */
  assign n5655_o = s_instr_category == 7'b1000100;
  /* control_fsm_rtl.vhd:1542:21  */
  assign n5657_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1545:24  */
  assign n5659_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1545:13  */
  assign n5662_o = n5659_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1545:13  */
  assign n5665_o = n5659_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1545:13  */
  assign n5668_o = n5659_o ? 4'b1111 : 4'b0000;
  /* control_fsm_rtl.vhd:1542:13  */
  assign n5671_o = n5657_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1542:13  */
  assign n5673_o = n5657_o ? 4'b0000 : n5662_o;
  /* control_fsm_rtl.vhd:1542:13  */
  assign n5675_o = n5657_o ? 3'b000 : n5665_o;
  /* control_fsm_rtl.vhd:1542:13  */
  assign n5677_o = n5657_o ? 4'b0000 : n5668_o;
  /* control_fsm_rtl.vhd:1542:13  */
  assign n5680_o = n5657_o ? 2'b01 : 2'b00;
  /* control_fsm_rtl.vhd:1541:11  */
  assign n5682_o = s_instr_category == 7'b1000101;
  /* control_fsm_rtl.vhd:1554:11  */
  assign n5684_o = s_instr_category == 7'b1000110;
  /* control_fsm_rtl.vhd:1562:11  */
  assign n5686_o = s_instr_category == 7'b1000111;
  /* control_fsm_rtl.vhd:1571:21  */
  assign n5688_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1574:24  */
  assign n5690_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1577:24  */
  assign n5692_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1577:13  */
  assign n5695_o = n5692_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1577:13  */
  assign n5698_o = n5692_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:1577:13  */
  assign n5701_o = n5692_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:1574:13  */
  assign n5704_o = n5690_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1574:13  */
  assign n5706_o = n5690_o ? 4'b0000 : n5695_o;
  /* control_fsm_rtl.vhd:1574:13  */
  assign n5708_o = n5690_o ? 3'b000 : n5698_o;
  /* control_fsm_rtl.vhd:1574:13  */
  assign n5710_o = n5690_o ? 4'b0000 : n5701_o;
  /* control_fsm_rtl.vhd:1574:13  */
  assign n5713_o = n5690_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1571:13  */
  assign n5715_o = n5688_o ? 3'b010 : n5704_o;
  /* control_fsm_rtl.vhd:1571:13  */
  assign n5717_o = n5688_o ? 4'b0001 : n5706_o;
  /* control_fsm_rtl.vhd:1571:13  */
  assign n5719_o = n5688_o ? 3'b000 : n5708_o;
  /* control_fsm_rtl.vhd:1571:13  */
  assign n5721_o = n5688_o ? 4'b0000 : n5710_o;
  /* control_fsm_rtl.vhd:1571:13  */
  assign n5723_o = n5688_o ? 4'b0000 : n5713_o;
  /* control_fsm_rtl.vhd:1570:11  */
  assign n5725_o = s_instr_category == 7'b1001000;
  /* control_fsm_rtl.vhd:1587:21  */
  assign n5727_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1590:24  */
  assign n5729_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1590:13  */
  assign n5732_o = n5729_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1590:13  */
  assign n5735_o = n5729_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:1590:13  */
  assign n5738_o = n5729_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1590:13  */
  assign n5741_o = n5729_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1587:13  */
  assign n5744_o = n5727_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1587:13  */
  assign n5746_o = n5727_o ? 4'b0001 : n5732_o;
  /* control_fsm_rtl.vhd:1587:13  */
  assign n5748_o = n5727_o ? 3'b000 : n5735_o;
  /* control_fsm_rtl.vhd:1587:13  */
  assign n5750_o = n5727_o ? 4'b0000 : n5738_o;
  /* control_fsm_rtl.vhd:1587:13  */
  assign n5752_o = n5727_o ? 4'b0000 : n5741_o;
  /* control_fsm_rtl.vhd:1586:11  */
  assign n5754_o = s_instr_category == 7'b1001001;
  /* control_fsm_rtl.vhd:1601:21  */
  assign n5756_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1604:24  */
  assign n5758_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1610:24  */
  assign n5760_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1610:13  */
  assign n5763_o = n5760_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1610:13  */
  assign n5766_o = n5760_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1610:13  */
  assign n5769_o = n5760_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:1610:13  */
  assign n5772_o = n5760_o ? 4'b1101 : 4'b0000;
  /* control_fsm_rtl.vhd:1604:13  */
  assign n5775_o = n5758_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1604:13  */
  assign n5777_o = n5758_o ? 4'b0001 : n5763_o;
  /* control_fsm_rtl.vhd:1604:13  */
  assign n5779_o = n5758_o ? 3'b100 : n5766_o;
  /* control_fsm_rtl.vhd:1604:13  */
  assign n5781_o = n5758_o ? 4'b0101 : n5769_o;
  /* control_fsm_rtl.vhd:1604:13  */
  assign n5783_o = n5758_o ? 4'b1110 : n5772_o;
  /* control_fsm_rtl.vhd:1601:13  */
  assign n5785_o = n5756_o ? 3'b010 : n5775_o;
  /* control_fsm_rtl.vhd:1601:13  */
  assign n5787_o = n5756_o ? 4'b0001 : n5777_o;
  /* control_fsm_rtl.vhd:1601:13  */
  assign n5789_o = n5756_o ? 3'b000 : n5779_o;
  /* control_fsm_rtl.vhd:1601:13  */
  assign n5791_o = n5756_o ? 4'b0000 : n5781_o;
  /* control_fsm_rtl.vhd:1601:13  */
  assign n5793_o = n5756_o ? 4'b0000 : n5783_o;
  /* control_fsm_rtl.vhd:1600:11  */
  assign n5795_o = s_instr_category == 7'b1001010;
  /* control_fsm_rtl.vhd:1621:21  */
  assign n5797_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1625:24  */
  assign n5799_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1630:24  */
  assign n5801_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1630:13  */
  assign n5804_o = n5801_o ? 6'b101010 : 6'b000000;
  /* control_fsm_rtl.vhd:1630:13  */
  assign n5807_o = n5801_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1630:13  */
  assign n5810_o = n5801_o ? 3'b111 : 3'b000;
  /* control_fsm_rtl.vhd:1630:13  */
  assign n5813_o = n5801_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1630:13  */
  assign n5816_o = n5801_o ? 4'b1100 : 4'b0000;
  /* control_fsm_rtl.vhd:1625:13  */
  assign n5818_o = n5799_o ? 6'b101010 : n5804_o;
  /* control_fsm_rtl.vhd:1625:13  */
  assign n5821_o = n5799_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1625:13  */
  assign n5823_o = n5799_o ? 4'b0000 : n5807_o;
  /* control_fsm_rtl.vhd:1625:13  */
  assign n5825_o = n5799_o ? 3'b000 : n5810_o;
  /* control_fsm_rtl.vhd:1625:13  */
  assign n5827_o = n5799_o ? 4'b0011 : n5813_o;
  /* control_fsm_rtl.vhd:1625:13  */
  assign n5829_o = n5799_o ? 4'b1100 : n5816_o;
  /* control_fsm_rtl.vhd:1621:13  */
  assign n5831_o = n5797_o ? 6'b101010 : n5818_o;
  /* control_fsm_rtl.vhd:1621:13  */
  assign n5833_o = n5797_o ? 3'b010 : n5821_o;
  /* control_fsm_rtl.vhd:1621:13  */
  assign n5835_o = n5797_o ? 4'b0000 : n5823_o;
  /* control_fsm_rtl.vhd:1621:13  */
  assign n5837_o = n5797_o ? 3'b000 : n5825_o;
  /* control_fsm_rtl.vhd:1621:13  */
  assign n5839_o = n5797_o ? 4'b0000 : n5827_o;
  /* control_fsm_rtl.vhd:1621:13  */
  assign n5841_o = n5797_o ? 4'b1100 : n5829_o;
  /* control_fsm_rtl.vhd:1620:11  */
  assign n5843_o = s_instr_category == 7'b1001011;
  /* control_fsm_rtl.vhd:1641:11  */
  assign n5845_o = s_instr_category == 7'b1001100;
  /* control_fsm_rtl.vhd:1648:21  */
  assign n5847_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1651:24  */
  assign n5849_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1651:13  */
  assign n5852_o = n5849_o ? 6'b101100 : 6'b000000;
  /* control_fsm_rtl.vhd:1651:13  */
  assign n5855_o = n5849_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1651:13  */
  assign n5858_o = n5849_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1651:13  */
  assign n5861_o = n5849_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1648:13  */
  assign n5863_o = n5847_o ? 6'b000000 : n5852_o;
  /* control_fsm_rtl.vhd:1648:13  */
  assign n5866_o = n5847_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1648:13  */
  assign n5868_o = n5847_o ? 4'b0000 : n5855_o;
  /* control_fsm_rtl.vhd:1648:13  */
  assign n5870_o = n5847_o ? 3'b000 : n5858_o;
  /* control_fsm_rtl.vhd:1648:13  */
  assign n5872_o = n5847_o ? 4'b0000 : n5861_o;
  /* control_fsm_rtl.vhd:1648:13  */
  assign n5875_o = n5847_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:1647:11  */
  assign n5877_o = s_instr_category == 7'b1001101;
  /* control_fsm_rtl.vhd:1661:21  */
  assign n5879_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1664:24  */
  assign n5881_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1667:24  */
  assign n5883_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1667:13  */
  assign n5886_o = n5883_o ? 6'b101100 : 6'b000000;
  /* control_fsm_rtl.vhd:1667:13  */
  assign n5889_o = n5883_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1667:13  */
  assign n5892_o = n5883_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1667:13  */
  assign n5895_o = n5883_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1664:13  */
  assign n5897_o = n5881_o ? 6'b000000 : n5886_o;
  /* control_fsm_rtl.vhd:1664:13  */
  assign n5900_o = n5881_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1664:13  */
  assign n5902_o = n5881_o ? 4'b0000 : n5889_o;
  /* control_fsm_rtl.vhd:1664:13  */
  assign n5904_o = n5881_o ? 3'b000 : n5892_o;
  /* control_fsm_rtl.vhd:1664:13  */
  assign n5906_o = n5881_o ? 4'b0000 : n5895_o;
  /* control_fsm_rtl.vhd:1664:13  */
  assign n5909_o = n5881_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1661:13  */
  assign n5911_o = n5879_o ? 6'b000000 : n5897_o;
  /* control_fsm_rtl.vhd:1661:13  */
  assign n5913_o = n5879_o ? 3'b010 : n5900_o;
  /* control_fsm_rtl.vhd:1661:13  */
  assign n5915_o = n5879_o ? 4'b0001 : n5902_o;
  /* control_fsm_rtl.vhd:1661:13  */
  assign n5917_o = n5879_o ? 3'b000 : n5904_o;
  /* control_fsm_rtl.vhd:1661:13  */
  assign n5919_o = n5879_o ? 4'b0000 : n5906_o;
  /* control_fsm_rtl.vhd:1661:13  */
  assign n5921_o = n5879_o ? 4'b0000 : n5909_o;
  /* control_fsm_rtl.vhd:1660:11  */
  assign n5923_o = s_instr_category == 7'b1001110;
  /* control_fsm_rtl.vhd:1677:21  */
  assign n5925_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1680:24  */
  assign n5927_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1680:13  */
  assign n5930_o = n5927_o ? 6'b101100 : 6'b000000;
  /* control_fsm_rtl.vhd:1680:13  */
  assign n5933_o = n5927_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1680:13  */
  assign n5936_o = n5927_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1680:13  */
  assign n5939_o = n5927_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1677:13  */
  assign n5941_o = n5925_o ? 6'b000000 : n5930_o;
  /* control_fsm_rtl.vhd:1677:13  */
  assign n5944_o = n5925_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1677:13  */
  assign n5946_o = n5925_o ? 4'b0000 : n5933_o;
  /* control_fsm_rtl.vhd:1677:13  */
  assign n5948_o = n5925_o ? 3'b000 : n5936_o;
  /* control_fsm_rtl.vhd:1677:13  */
  assign n5950_o = n5925_o ? 4'b0000 : n5939_o;
  /* control_fsm_rtl.vhd:1677:13  */
  assign n5953_o = n5925_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:1676:11  */
  assign n5955_o = s_instr_category == 7'b1001111;
  /* control_fsm_rtl.vhd:1690:21  */
  assign n5957_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1693:24  */
  assign n5959_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1693:13  */
  assign n5962_o = n5959_o ? 6'b101101 : 6'b000000;
  /* control_fsm_rtl.vhd:1693:13  */
  assign n5965_o = n5959_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1693:13  */
  assign n5968_o = n5959_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:1693:13  */
  assign n5971_o = n5959_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1690:13  */
  assign n5973_o = n5957_o ? 6'b000000 : n5962_o;
  /* control_fsm_rtl.vhd:1690:13  */
  assign n5976_o = n5957_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1690:13  */
  assign n5978_o = n5957_o ? 4'b0001 : n5965_o;
  /* control_fsm_rtl.vhd:1690:13  */
  assign n5980_o = n5957_o ? 3'b000 : n5968_o;
  /* control_fsm_rtl.vhd:1690:13  */
  assign n5982_o = n5957_o ? 4'b0000 : n5971_o;
  /* control_fsm_rtl.vhd:1689:11  */
  assign n5984_o = s_instr_category == 7'b1010000;
  /* control_fsm_rtl.vhd:1703:21  */
  assign n5986_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1706:24  */
  assign n5988_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1709:24  */
  assign n5990_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1709:13  */
  assign n5993_o = n5990_o ? 6'b101100 : 6'b000000;
  /* control_fsm_rtl.vhd:1709:13  */
  assign n5996_o = n5990_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1709:13  */
  assign n5999_o = n5990_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1709:13  */
  assign n6002_o = n5990_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1709:13  */
  assign n6005_o = n5990_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1706:13  */
  assign n6007_o = n5988_o ? 6'b000000 : n5993_o;
  /* control_fsm_rtl.vhd:1706:13  */
  assign n6010_o = n5988_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1706:13  */
  assign n6012_o = n5988_o ? 4'b0000 : n5996_o;
  /* control_fsm_rtl.vhd:1706:13  */
  assign n6014_o = n5988_o ? 3'b000 : n5999_o;
  /* control_fsm_rtl.vhd:1706:13  */
  assign n6016_o = n5988_o ? 4'b0000 : n6002_o;
  /* control_fsm_rtl.vhd:1706:13  */
  assign n6018_o = n5988_o ? 4'b1000 : n6005_o;
  /* control_fsm_rtl.vhd:1703:13  */
  assign n6020_o = n5986_o ? 6'b000000 : n6007_o;
  /* control_fsm_rtl.vhd:1703:13  */
  assign n6022_o = n5986_o ? 3'b010 : n6010_o;
  /* control_fsm_rtl.vhd:1703:13  */
  assign n6024_o = n5986_o ? 4'b0001 : n6012_o;
  /* control_fsm_rtl.vhd:1703:13  */
  assign n6026_o = n5986_o ? 3'b000 : n6014_o;
  /* control_fsm_rtl.vhd:1703:13  */
  assign n6028_o = n5986_o ? 4'b0000 : n6016_o;
  /* control_fsm_rtl.vhd:1703:13  */
  assign n6030_o = n5986_o ? 4'b0000 : n6018_o;
  /* control_fsm_rtl.vhd:1702:11  */
  assign n6032_o = s_instr_category == 7'b1010001;
  /* control_fsm_rtl.vhd:1721:21  */
  assign n6034_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1724:24  */
  assign n6036_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1729:24  */
  assign n6038_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1729:13  */
  assign n6041_o = n6038_o ? 6'b101110 : 6'b000000;
  /* control_fsm_rtl.vhd:1729:13  */
  assign n6044_o = n6038_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1729:13  */
  assign n6047_o = n6038_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1729:13  */
  assign n6050_o = n6038_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1729:13  */
  assign n6053_o = n6038_o ? 4'b1010 : 4'b0000;
  /* control_fsm_rtl.vhd:1724:13  */
  assign n6055_o = n6036_o ? 6'b000000 : n6041_o;
  /* control_fsm_rtl.vhd:1724:13  */
  assign n6058_o = n6036_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1724:13  */
  assign n6060_o = n6036_o ? 4'b0001 : n6044_o;
  /* control_fsm_rtl.vhd:1724:13  */
  assign n6062_o = n6036_o ? 3'b000 : n6047_o;
  /* control_fsm_rtl.vhd:1724:13  */
  assign n6064_o = n6036_o ? 4'b0000 : n6050_o;
  /* control_fsm_rtl.vhd:1724:13  */
  assign n6066_o = n6036_o ? 4'b1000 : n6053_o;
  /* control_fsm_rtl.vhd:1724:13  */
  assign n6069_o = n6036_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1721:13  */
  assign n6071_o = n6034_o ? 6'b000000 : n6055_o;
  /* control_fsm_rtl.vhd:1721:13  */
  assign n6073_o = n6034_o ? 3'b010 : n6058_o;
  /* control_fsm_rtl.vhd:1721:13  */
  assign n6075_o = n6034_o ? 4'b0001 : n6060_o;
  /* control_fsm_rtl.vhd:1721:13  */
  assign n6077_o = n6034_o ? 3'b000 : n6062_o;
  /* control_fsm_rtl.vhd:1721:13  */
  assign n6079_o = n6034_o ? 4'b0000 : n6064_o;
  /* control_fsm_rtl.vhd:1721:13  */
  assign n6081_o = n6034_o ? 4'b0000 : n6066_o;
  /* control_fsm_rtl.vhd:1721:13  */
  assign n6083_o = n6034_o ? 4'b0000 : n6069_o;
  /* control_fsm_rtl.vhd:1720:11  */
  assign n6085_o = s_instr_category == 7'b1010010;
  /* control_fsm_rtl.vhd:1741:21  */
  assign n6087_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1744:24  */
  assign n6089_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1747:24  */
  assign n6091_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1747:13  */
  assign n6094_o = n6091_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1747:13  */
  assign n6097_o = n6091_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:1747:13  */
  assign n6100_o = n6091_o ? 4'b1001 : 4'b0000;
  /* control_fsm_rtl.vhd:1744:13  */
  assign n6103_o = n6089_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1744:13  */
  assign n6105_o = n6089_o ? 4'b0000 : n6094_o;
  /* control_fsm_rtl.vhd:1744:13  */
  assign n6107_o = n6089_o ? 3'b000 : n6097_o;
  /* control_fsm_rtl.vhd:1744:13  */
  assign n6109_o = n6089_o ? 4'b0000 : n6100_o;
  /* control_fsm_rtl.vhd:1744:13  */
  assign n6112_o = n6089_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1741:13  */
  assign n6114_o = n6087_o ? 3'b010 : n6103_o;
  /* control_fsm_rtl.vhd:1741:13  */
  assign n6116_o = n6087_o ? 4'b0001 : n6105_o;
  /* control_fsm_rtl.vhd:1741:13  */
  assign n6118_o = n6087_o ? 3'b000 : n6107_o;
  /* control_fsm_rtl.vhd:1741:13  */
  assign n6120_o = n6087_o ? 4'b0000 : n6109_o;
  /* control_fsm_rtl.vhd:1741:13  */
  assign n6122_o = n6087_o ? 4'b0000 : n6112_o;
  /* control_fsm_rtl.vhd:1740:11  */
  assign n6124_o = s_instr_category == 7'b1010011;
  /* control_fsm_rtl.vhd:1757:21  */
  assign n6126_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1760:24  */
  assign n6128_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1763:24  */
  assign n6130_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1763:13  */
  assign n6133_o = n6130_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1763:13  */
  assign n6136_o = n6130_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:1763:13  */
  assign n6139_o = n6130_o ? 4'b1010 : 4'b0000;
  /* control_fsm_rtl.vhd:1760:13  */
  assign n6142_o = n6128_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1760:13  */
  assign n6144_o = n6128_o ? 4'b0000 : n6133_o;
  /* control_fsm_rtl.vhd:1760:13  */
  assign n6146_o = n6128_o ? 3'b000 : n6136_o;
  /* control_fsm_rtl.vhd:1760:13  */
  assign n6148_o = n6128_o ? 4'b0000 : n6139_o;
  /* control_fsm_rtl.vhd:1760:13  */
  assign n6151_o = n6128_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1757:13  */
  assign n6153_o = n6126_o ? 3'b010 : n6142_o;
  /* control_fsm_rtl.vhd:1757:13  */
  assign n6155_o = n6126_o ? 4'b0001 : n6144_o;
  /* control_fsm_rtl.vhd:1757:13  */
  assign n6157_o = n6126_o ? 3'b000 : n6146_o;
  /* control_fsm_rtl.vhd:1757:13  */
  assign n6159_o = n6126_o ? 4'b0000 : n6148_o;
  /* control_fsm_rtl.vhd:1757:13  */
  assign n6161_o = n6126_o ? 4'b0000 : n6151_o;
  /* control_fsm_rtl.vhd:1756:11  */
  assign n6163_o = s_instr_category == 7'b1010100;
  /* control_fsm_rtl.vhd:1773:21  */
  assign n6165_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1777:24  */
  assign n6167_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1777:13  */
  assign n6170_o = n6167_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1777:13  */
  assign n6173_o = n6167_o ? 3'b101 : 3'b000;
  /* control_fsm_rtl.vhd:1777:13  */
  assign n6176_o = n6167_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1777:13  */
  assign n6179_o = n6167_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1773:13  */
  assign n6182_o = n6165_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1773:13  */
  assign n6184_o = n6165_o ? 4'b0001 : n6170_o;
  /* control_fsm_rtl.vhd:1773:13  */
  assign n6186_o = n6165_o ? 3'b000 : n6173_o;
  /* control_fsm_rtl.vhd:1773:13  */
  assign n6188_o = n6165_o ? 4'b0000 : n6176_o;
  /* control_fsm_rtl.vhd:1773:13  */
  assign n6190_o = n6165_o ? 4'b0101 : n6179_o;
  /* control_fsm_rtl.vhd:1772:11  */
  assign n6192_o = s_instr_category == 7'b1010101;
  /* control_fsm_rtl.vhd:1788:21  */
  assign n6194_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1792:24  */
  assign n6196_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1795:24  */
  assign n6198_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1795:13  */
  assign n6201_o = n6198_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1795:13  */
  assign n6204_o = n6198_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:1795:13  */
  assign n6207_o = n6198_o ? 4'b0100 : 4'b0000;
  /* control_fsm_rtl.vhd:1795:13  */
  assign n6210_o = n6198_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:1792:13  */
  assign n6213_o = n6196_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1792:13  */
  assign n6215_o = n6196_o ? 4'b0000 : n6201_o;
  /* control_fsm_rtl.vhd:1792:13  */
  assign n6217_o = n6196_o ? 3'b000 : n6204_o;
  /* control_fsm_rtl.vhd:1792:13  */
  assign n6219_o = n6196_o ? 4'b0000 : n6207_o;
  /* control_fsm_rtl.vhd:1792:13  */
  assign n6221_o = n6196_o ? 4'b1000 : n6210_o;
  /* control_fsm_rtl.vhd:1788:13  */
  assign n6223_o = n6194_o ? 3'b010 : n6213_o;
  /* control_fsm_rtl.vhd:1788:13  */
  assign n6225_o = n6194_o ? 4'b0001 : n6215_o;
  /* control_fsm_rtl.vhd:1788:13  */
  assign n6227_o = n6194_o ? 3'b001 : n6217_o;
  /* control_fsm_rtl.vhd:1788:13  */
  assign n6229_o = n6194_o ? 4'b0000 : n6219_o;
  /* control_fsm_rtl.vhd:1788:13  */
  assign n6231_o = n6194_o ? 4'b0000 : n6221_o;
  /* control_fsm_rtl.vhd:1787:11  */
  assign n6233_o = s_instr_category == 7'b1010110;
  /* control_fsm_rtl.vhd:1806:21  */
  assign n6235_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1810:24  */
  assign n6237_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1814:24  */
  assign n6239_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1814:13  */
  assign n6242_o = n6239_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1814:13  */
  assign n6245_o = n6239_o ? 3'b001 : 3'b000;
  /* control_fsm_rtl.vhd:1810:13  */
  assign n6248_o = n6237_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1810:13  */
  assign n6250_o = n6237_o ? 4'b0000 : n6242_o;
  /* control_fsm_rtl.vhd:1810:13  */
  assign n6252_o = n6237_o ? 3'b000 : n6245_o;
  /* control_fsm_rtl.vhd:1810:13  */
  assign n6255_o = n6237_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:1810:13  */
  assign n6258_o = n6237_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1806:13  */
  assign n6260_o = n6235_o ? 3'b010 : n6248_o;
  /* control_fsm_rtl.vhd:1806:13  */
  assign n6262_o = n6235_o ? 4'b0000 : n6250_o;
  /* control_fsm_rtl.vhd:1806:13  */
  assign n6264_o = n6235_o ? 3'b001 : n6252_o;
  /* control_fsm_rtl.vhd:1806:13  */
  assign n6266_o = n6235_o ? 4'b0101 : n6255_o;
  /* control_fsm_rtl.vhd:1806:13  */
  assign n6268_o = n6235_o ? 4'b0000 : n6258_o;
  /* control_fsm_rtl.vhd:1805:11  */
  assign n6270_o = s_instr_category == 7'b1010111;
  /* control_fsm_rtl.vhd:1823:21  */
  assign n6272_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1827:24  */
  assign n6274_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1831:24  */
  assign n6276_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1839:15  */
  assign n6279_o = s_intlow ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:1839:15  */
  assign n6282_o = s_intlow ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:1839:15  */
  assign n6285_o = s_intlow ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:1832:15  */
  assign n6287_o = s_inthigh ? 1'b0 : n6279_o;
  /* control_fsm_rtl.vhd:1832:15  */
  assign n6290_o = s_inthigh ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:1832:15  */
  assign n6292_o = s_inthigh ? 1'b0 : n6282_o;
  /* control_fsm_rtl.vhd:1832:15  */
  assign n6294_o = s_inthigh ? 1'b0 : n6285_o;
  /* control_fsm_rtl.vhd:1832:15  */
  assign n6297_o = s_inthigh ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:1832:15  */
  assign n6300_o = s_inthigh ? 1'b1 : 1'b0;
  /* control_fsm_rtl.vhd:1831:13  */
  assign n6303_o = n6276_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1831:13  */
  assign n6306_o = n6276_o ? 3'b001 : 3'b000;
  /* control_fsm_rtl.vhd:1831:13  */
  assign n6308_o = n6276_o ? n6287_o : 1'b0;
  /* control_fsm_rtl.vhd:1831:13  */
  assign n6310_o = n6276_o ? n6290_o : 1'b0;
  /* control_fsm_rtl.vhd:1831:13  */
  assign n6312_o = n6276_o ? n6292_o : 1'b0;
  /* control_fsm_rtl.vhd:1831:13  */
  assign n6314_o = n6276_o ? n6294_o : 1'b0;
  /* control_fsm_rtl.vhd:1831:13  */
  assign n6316_o = n6276_o ? n6297_o : 1'b0;
  /* control_fsm_rtl.vhd:1831:13  */
  assign n6318_o = n6276_o ? n6300_o : 1'b0;
  /* control_fsm_rtl.vhd:1827:13  */
  assign n6321_o = n6274_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1827:13  */
  assign n6323_o = n6274_o ? 4'b0000 : n6303_o;
  /* control_fsm_rtl.vhd:1827:13  */
  assign n6325_o = n6274_o ? 3'b000 : n6306_o;
  /* control_fsm_rtl.vhd:1827:13  */
  assign n6328_o = n6274_o ? 4'b0101 : 4'b0000;
  /* control_fsm_rtl.vhd:1827:13  */
  assign n6331_o = n6274_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1827:13  */
  assign n6333_o = n6274_o ? 1'b0 : n6308_o;
  /* control_fsm_rtl.vhd:1827:13  */
  assign n6335_o = n6274_o ? 1'b0 : n6310_o;
  /* control_fsm_rtl.vhd:1827:13  */
  assign n6337_o = n6274_o ? 1'b0 : n6312_o;
  /* control_fsm_rtl.vhd:1827:13  */
  assign n6339_o = n6274_o ? 1'b0 : n6314_o;
  /* control_fsm_rtl.vhd:1827:13  */
  assign n6341_o = n6274_o ? 1'b0 : n6316_o;
  /* control_fsm_rtl.vhd:1827:13  */
  assign n6343_o = n6274_o ? 1'b0 : n6318_o;
  /* control_fsm_rtl.vhd:1823:13  */
  assign n6345_o = n6272_o ? 3'b010 : n6321_o;
  /* control_fsm_rtl.vhd:1823:13  */
  assign n6347_o = n6272_o ? 4'b0000 : n6323_o;
  /* control_fsm_rtl.vhd:1823:13  */
  assign n6349_o = n6272_o ? 3'b001 : n6325_o;
  /* control_fsm_rtl.vhd:1823:13  */
  assign n6351_o = n6272_o ? 4'b0101 : n6328_o;
  /* control_fsm_rtl.vhd:1823:13  */
  assign n6353_o = n6272_o ? 4'b0000 : n6331_o;
  /* control_fsm_rtl.vhd:1823:13  */
  assign n6355_o = n6272_o ? 1'b0 : n6333_o;
  /* control_fsm_rtl.vhd:1823:13  */
  assign n6357_o = n6272_o ? 1'b0 : n6335_o;
  /* control_fsm_rtl.vhd:1823:13  */
  assign n6359_o = n6272_o ? 1'b0 : n6337_o;
  /* control_fsm_rtl.vhd:1823:13  */
  assign n6361_o = n6272_o ? 1'b0 : n6339_o;
  /* control_fsm_rtl.vhd:1823:13  */
  assign n6363_o = n6272_o ? 1'b0 : n6341_o;
  /* control_fsm_rtl.vhd:1823:13  */
  assign n6365_o = n6272_o ? 1'b0 : n6343_o;
  /* control_fsm_rtl.vhd:1822:11  */
  assign n6367_o = s_instr_category == 7'b1011000;
  /* control_fsm_rtl.vhd:1856:11  */
  assign n6369_o = s_instr_category == 7'b1011001;
  /* control_fsm_rtl.vhd:1865:11  */
  assign n6371_o = s_instr_category == 7'b1011010;
  /* control_fsm_rtl.vhd:1874:11  */
  assign n6373_o = s_instr_category == 7'b1011011;
  /* control_fsm_rtl.vhd:1883:11  */
  assign n6375_o = s_instr_category == 7'b1011100;
  /* control_fsm_rtl.vhd:1892:11  */
  assign n6377_o = s_instr_category == 7'b1011101;
  /* control_fsm_rtl.vhd:1902:21  */
  assign n6379_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1905:24  */
  assign n6381_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1905:13  */
  assign n6384_o = n6381_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1905:13  */
  assign n6387_o = n6381_o ? 3'b110 : 3'b000;
  /* control_fsm_rtl.vhd:1905:13  */
  assign n6390_o = n6381_o ? 4'b1011 : 4'b0000;
  /* control_fsm_rtl.vhd:1905:13  */
  assign n6393_o = n6381_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1902:13  */
  assign n6396_o = n6379_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1902:13  */
  assign n6398_o = n6379_o ? 4'b0001 : n6384_o;
  /* control_fsm_rtl.vhd:1902:13  */
  assign n6400_o = n6379_o ? 3'b000 : n6387_o;
  /* control_fsm_rtl.vhd:1902:13  */
  assign n6402_o = n6379_o ? 4'b0000 : n6390_o;
  /* control_fsm_rtl.vhd:1902:13  */
  assign n6404_o = n6379_o ? 4'b0000 : n6393_o;
  /* control_fsm_rtl.vhd:1901:11  */
  assign n6406_o = s_instr_category == 7'b1011110;
  /* control_fsm_rtl.vhd:1916:21  */
  assign n6408_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1919:24  */
  assign n6410_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1919:13  */
  assign n6413_o = n6410_o ? 4'b0010 : 4'b0000;
  /* control_fsm_rtl.vhd:1916:13  */
  assign n6416_o = n6408_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1916:13  */
  assign n6418_o = n6408_o ? 4'b0001 : n6413_o;
  /* control_fsm_rtl.vhd:1915:11  */
  assign n6420_o = s_instr_category == 7'b1011111;
  /* control_fsm_rtl.vhd:1927:21  */
  assign n6422_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1930:24  */
  assign n6424_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1930:13  */
  assign n6427_o = n6424_o ? 6'b101000 : 6'b000000;
  /* control_fsm_rtl.vhd:1930:13  */
  assign n6430_o = n6424_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1930:13  */
  assign n6433_o = n6424_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:1930:13  */
  assign n6436_o = n6424_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1927:13  */
  assign n6438_o = n6422_o ? 6'b000000 : n6427_o;
  /* control_fsm_rtl.vhd:1927:13  */
  assign n6441_o = n6422_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1927:13  */
  assign n6443_o = n6422_o ? 4'b0000 : n6430_o;
  /* control_fsm_rtl.vhd:1927:13  */
  assign n6445_o = n6422_o ? 3'b000 : n6433_o;
  /* control_fsm_rtl.vhd:1927:13  */
  assign n6447_o = n6422_o ? 4'b0000 : n6436_o;
  /* control_fsm_rtl.vhd:1927:13  */
  assign n6450_o = n6422_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:1926:11  */
  assign n6452_o = s_instr_category == 7'b1100000;
  /* control_fsm_rtl.vhd:1940:21  */
  assign n6454_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1943:24  */
  assign n6456_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1946:24  */
  assign n6458_o = state == 3'b011;
  /* control_fsm_rtl.vhd:1946:13  */
  assign n6461_o = n6458_o ? 6'b101000 : 6'b000000;
  /* control_fsm_rtl.vhd:1946:13  */
  assign n6464_o = n6458_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1946:13  */
  assign n6467_o = n6458_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:1946:13  */
  assign n6470_o = n6458_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1943:13  */
  assign n6472_o = n6456_o ? 6'b000000 : n6461_o;
  /* control_fsm_rtl.vhd:1943:13  */
  assign n6475_o = n6456_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1943:13  */
  assign n6477_o = n6456_o ? 4'b0000 : n6464_o;
  /* control_fsm_rtl.vhd:1943:13  */
  assign n6479_o = n6456_o ? 3'b000 : n6467_o;
  /* control_fsm_rtl.vhd:1943:13  */
  assign n6481_o = n6456_o ? 4'b0000 : n6470_o;
  /* control_fsm_rtl.vhd:1943:13  */
  assign n6484_o = n6456_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1940:13  */
  assign n6486_o = n6454_o ? 6'b000000 : n6472_o;
  /* control_fsm_rtl.vhd:1940:13  */
  assign n6488_o = n6454_o ? 3'b010 : n6475_o;
  /* control_fsm_rtl.vhd:1940:13  */
  assign n6490_o = n6454_o ? 4'b0001 : n6477_o;
  /* control_fsm_rtl.vhd:1940:13  */
  assign n6492_o = n6454_o ? 3'b000 : n6479_o;
  /* control_fsm_rtl.vhd:1940:13  */
  assign n6494_o = n6454_o ? 4'b0000 : n6481_o;
  /* control_fsm_rtl.vhd:1940:13  */
  assign n6496_o = n6454_o ? 4'b0000 : n6484_o;
  /* control_fsm_rtl.vhd:1939:11  */
  assign n6498_o = s_instr_category == 7'b1100001;
  /* control_fsm_rtl.vhd:1956:21  */
  assign n6500_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1959:24  */
  assign n6502_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1959:13  */
  assign n6505_o = n6502_o ? 6'b101000 : 6'b000000;
  /* control_fsm_rtl.vhd:1959:13  */
  assign n6508_o = n6502_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1959:13  */
  assign n6511_o = n6502_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:1959:13  */
  assign n6514_o = n6502_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1956:13  */
  assign n6516_o = n6500_o ? 6'b000000 : n6505_o;
  /* control_fsm_rtl.vhd:1956:13  */
  assign n6519_o = n6500_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1956:13  */
  assign n6521_o = n6500_o ? 4'b0000 : n6508_o;
  /* control_fsm_rtl.vhd:1956:13  */
  assign n6523_o = n6500_o ? 3'b000 : n6511_o;
  /* control_fsm_rtl.vhd:1956:13  */
  assign n6525_o = n6500_o ? 4'b0000 : n6514_o;
  /* control_fsm_rtl.vhd:1956:13  */
  assign n6528_o = n6500_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:1955:11  */
  assign n6530_o = s_instr_category == 7'b1100010;
  /* control_fsm_rtl.vhd:1970:21  */
  assign n6532_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1973:24  */
  assign n6534_o = state == 3'b010;
  /* control_fsm_rtl.vhd:1973:13  */
  assign n6537_o = n6534_o ? 6'b101001 : 6'b000000;
  /* control_fsm_rtl.vhd:1973:13  */
  assign n6540_o = n6534_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:1973:13  */
  assign n6543_o = n6534_o ? 3'b011 : 3'b000;
  /* control_fsm_rtl.vhd:1973:13  */
  assign n6546_o = n6534_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1970:13  */
  assign n6548_o = n6532_o ? 6'b000000 : n6537_o;
  /* control_fsm_rtl.vhd:1970:13  */
  assign n6551_o = n6532_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:1970:13  */
  assign n6553_o = n6532_o ? 4'b0001 : n6540_o;
  /* control_fsm_rtl.vhd:1970:13  */
  assign n6555_o = n6532_o ? 3'b000 : n6543_o;
  /* control_fsm_rtl.vhd:1970:13  */
  assign n6557_o = n6532_o ? 4'b0000 : n6546_o;
  /* control_fsm_rtl.vhd:1969:11  */
  assign n6559_o = s_instr_category == 7'b1100011;
  /* control_fsm_rtl.vhd:1983:11  */
  assign n6561_o = s_instr_category == 7'b1100100;
  /* control_fsm_rtl.vhd:1992:21  */
  assign n6563_o = state == 3'b001;
  /* control_fsm_rtl.vhd:1995:24  */
  assign n6565_o = state == 3'b010;
  /* control_fsm_rtl.vhd:2001:24  */
  assign n6567_o = state == 3'b011;
  /* control_fsm_rtl.vhd:2001:13  */
  assign n6570_o = n6567_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:2001:13  */
  assign n6573_o = n6567_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:2001:13  */
  assign n6576_o = n6567_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:1995:13  */
  assign n6579_o = n6565_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:1995:13  */
  assign n6581_o = n6565_o ? 4'b0000 : n6570_o;
  /* control_fsm_rtl.vhd:1995:13  */
  assign n6583_o = n6565_o ? 3'b100 : n6573_o;
  /* control_fsm_rtl.vhd:1995:13  */
  assign n6585_o = n6565_o ? 4'b0110 : n6576_o;
  /* control_fsm_rtl.vhd:1995:13  */
  assign n6588_o = n6565_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:1995:13  */
  assign n6591_o = n6565_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:1992:13  */
  assign n6593_o = n6563_o ? 3'b010 : n6579_o;
  /* control_fsm_rtl.vhd:1992:13  */
  assign n6595_o = n6563_o ? 4'b0000 : n6581_o;
  /* control_fsm_rtl.vhd:1992:13  */
  assign n6597_o = n6563_o ? 3'b000 : n6583_o;
  /* control_fsm_rtl.vhd:1992:13  */
  assign n6599_o = n6563_o ? 4'b0000 : n6585_o;
  /* control_fsm_rtl.vhd:1992:13  */
  assign n6601_o = n6563_o ? 4'b0110 : n6588_o;
  /* control_fsm_rtl.vhd:1992:13  */
  assign n6603_o = n6563_o ? 4'b0000 : n6591_o;
  /* control_fsm_rtl.vhd:1991:11  */
  assign n6605_o = s_instr_category == 7'b1100101;
  /* control_fsm_rtl.vhd:2011:21  */
  assign n6607_o = state == 3'b001;
  /* control_fsm_rtl.vhd:2014:24  */
  assign n6609_o = state == 3'b010;
  /* control_fsm_rtl.vhd:2017:24  */
  assign n6611_o = state == 3'b011;
  /* control_fsm_rtl.vhd:2023:24  */
  assign n6613_o = state == 3'b100;
  /* control_fsm_rtl.vhd:2023:13  */
  assign n6616_o = n6613_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:2023:13  */
  assign n6619_o = n6613_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:2023:13  */
  assign n6622_o = n6613_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:2017:13  */
  assign n6625_o = n6611_o ? 3'b100 : 3'b001;
  /* control_fsm_rtl.vhd:2017:13  */
  assign n6627_o = n6611_o ? 4'b0000 : n6616_o;
  /* control_fsm_rtl.vhd:2017:13  */
  assign n6629_o = n6611_o ? 3'b100 : n6619_o;
  /* control_fsm_rtl.vhd:2017:13  */
  assign n6631_o = n6611_o ? 4'b0110 : n6622_o;
  /* control_fsm_rtl.vhd:2017:13  */
  assign n6634_o = n6611_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:2017:13  */
  assign n6637_o = n6611_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:2014:13  */
  assign n6639_o = n6609_o ? 3'b011 : n6625_o;
  /* control_fsm_rtl.vhd:2014:13  */
  assign n6641_o = n6609_o ? 4'b0000 : n6627_o;
  /* control_fsm_rtl.vhd:2014:13  */
  assign n6643_o = n6609_o ? 3'b000 : n6629_o;
  /* control_fsm_rtl.vhd:2014:13  */
  assign n6645_o = n6609_o ? 4'b0000 : n6631_o;
  /* control_fsm_rtl.vhd:2014:13  */
  assign n6647_o = n6609_o ? 4'b1000 : n6634_o;
  /* control_fsm_rtl.vhd:2014:13  */
  assign n6649_o = n6609_o ? 4'b0000 : n6637_o;
  /* control_fsm_rtl.vhd:2011:13  */
  assign n6651_o = n6607_o ? 3'b010 : n6639_o;
  /* control_fsm_rtl.vhd:2011:13  */
  assign n6653_o = n6607_o ? 4'b0001 : n6641_o;
  /* control_fsm_rtl.vhd:2011:13  */
  assign n6655_o = n6607_o ? 3'b000 : n6643_o;
  /* control_fsm_rtl.vhd:2011:13  */
  assign n6657_o = n6607_o ? 4'b0000 : n6645_o;
  /* control_fsm_rtl.vhd:2011:13  */
  assign n6659_o = n6607_o ? 4'b0000 : n6647_o;
  /* control_fsm_rtl.vhd:2011:13  */
  assign n6661_o = n6607_o ? 4'b0000 : n6649_o;
  /* control_fsm_rtl.vhd:2010:11  */
  assign n6663_o = s_instr_category == 7'b1100110;
  /* control_fsm_rtl.vhd:2033:21  */
  assign n6665_o = state == 3'b001;
  /* control_fsm_rtl.vhd:2036:24  */
  assign n6667_o = state == 3'b010;
  /* control_fsm_rtl.vhd:2042:24  */
  assign n6669_o = state == 3'b011;
  /* control_fsm_rtl.vhd:2042:13  */
  assign n6672_o = n6669_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:2042:13  */
  assign n6675_o = n6669_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:2042:13  */
  assign n6678_o = n6669_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:2036:13  */
  assign n6681_o = n6667_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:2036:13  */
  assign n6683_o = n6667_o ? 4'b0000 : n6672_o;
  /* control_fsm_rtl.vhd:2036:13  */
  assign n6685_o = n6667_o ? 3'b100 : n6675_o;
  /* control_fsm_rtl.vhd:2036:13  */
  assign n6687_o = n6667_o ? 4'b0110 : n6678_o;
  /* control_fsm_rtl.vhd:2036:13  */
  assign n6690_o = n6667_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:2036:13  */
  assign n6693_o = n6667_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:2033:13  */
  assign n6695_o = n6665_o ? 3'b010 : n6681_o;
  /* control_fsm_rtl.vhd:2033:13  */
  assign n6697_o = n6665_o ? 4'b0000 : n6683_o;
  /* control_fsm_rtl.vhd:2033:13  */
  assign n6699_o = n6665_o ? 3'b000 : n6685_o;
  /* control_fsm_rtl.vhd:2033:13  */
  assign n6701_o = n6665_o ? 4'b0000 : n6687_o;
  /* control_fsm_rtl.vhd:2033:13  */
  assign n6703_o = n6665_o ? 4'b0111 : n6690_o;
  /* control_fsm_rtl.vhd:2033:13  */
  assign n6705_o = n6665_o ? 4'b0000 : n6693_o;
  /* control_fsm_rtl.vhd:2032:11  */
  assign n6707_o = s_instr_category == 7'b1100111;
  /* control_fsm_rtl.vhd:2052:21  */
  assign n6709_o = state == 3'b001;
  /* control_fsm_rtl.vhd:2056:24  */
  assign n6711_o = state == 3'b010;
  /* control_fsm_rtl.vhd:2061:24  */
  assign n6713_o = state == 3'b011;
  /* control_fsm_rtl.vhd:2061:13  */
  assign n6716_o = n6713_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:2061:13  */
  assign n6719_o = n6713_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:2061:13  */
  assign n6722_o = n6713_o ? 4'b1001 : 4'b0000;
  /* control_fsm_rtl.vhd:2061:13  */
  assign n6725_o = n6713_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:2056:13  */
  assign n6728_o = n6711_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:2056:13  */
  assign n6730_o = n6711_o ? 4'b0000 : n6716_o;
  /* control_fsm_rtl.vhd:2056:13  */
  assign n6732_o = n6711_o ? 3'b010 : n6719_o;
  /* control_fsm_rtl.vhd:2056:13  */
  assign n6734_o = n6711_o ? 4'b1010 : n6722_o;
  /* control_fsm_rtl.vhd:2056:13  */
  assign n6736_o = n6711_o ? 4'b0111 : n6725_o;
  /* control_fsm_rtl.vhd:2052:13  */
  assign n6738_o = n6709_o ? 3'b010 : n6728_o;
  /* control_fsm_rtl.vhd:2052:13  */
  assign n6740_o = n6709_o ? 4'b0000 : n6730_o;
  /* control_fsm_rtl.vhd:2052:13  */
  assign n6742_o = n6709_o ? 3'b000 : n6732_o;
  /* control_fsm_rtl.vhd:2052:13  */
  assign n6744_o = n6709_o ? 4'b0000 : n6734_o;
  /* control_fsm_rtl.vhd:2052:13  */
  assign n6746_o = n6709_o ? 4'b0111 : n6736_o;
  /* control_fsm_rtl.vhd:2052:13  */
  assign n6749_o = n6709_o ? 4'b1010 : 4'b0000;
  /* control_fsm_rtl.vhd:2051:11  */
  assign n6751_o = s_instr_category == 7'b1101000;
  /* control_fsm_rtl.vhd:2072:21  */
  assign n6753_o = state == 3'b001;
  /* control_fsm_rtl.vhd:2075:24  */
  assign n6755_o = state == 3'b010;
  /* control_fsm_rtl.vhd:2075:13  */
  assign n6758_o = n6755_o ? 6'b101111 : 6'b000000;
  /* control_fsm_rtl.vhd:2075:13  */
  assign n6761_o = n6755_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:2075:13  */
  assign n6764_o = n6755_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:2075:13  */
  assign n6767_o = n6755_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:2072:13  */
  assign n6769_o = n6753_o ? 6'b000000 : n6758_o;
  /* control_fsm_rtl.vhd:2072:13  */
  assign n6772_o = n6753_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:2072:13  */
  assign n6774_o = n6753_o ? 4'b0000 : n6761_o;
  /* control_fsm_rtl.vhd:2072:13  */
  assign n6776_o = n6753_o ? 3'b000 : n6764_o;
  /* control_fsm_rtl.vhd:2072:13  */
  assign n6778_o = n6753_o ? 4'b0000 : n6767_o;
  /* control_fsm_rtl.vhd:2072:13  */
  assign n6781_o = n6753_o ? 4'b0110 : 4'b0000;
  /* control_fsm_rtl.vhd:2071:11  */
  assign n6783_o = s_instr_category == 7'b1101001;
  /* control_fsm_rtl.vhd:2085:21  */
  assign n6785_o = state == 3'b001;
  /* control_fsm_rtl.vhd:2088:24  */
  assign n6787_o = state == 3'b010;
  /* control_fsm_rtl.vhd:2091:24  */
  assign n6789_o = state == 3'b011;
  /* control_fsm_rtl.vhd:2091:13  */
  assign n6792_o = n6789_o ? 6'b101111 : 6'b000000;
  /* control_fsm_rtl.vhd:2091:13  */
  assign n6795_o = n6789_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:2091:13  */
  assign n6798_o = n6789_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:2091:13  */
  assign n6801_o = n6789_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:2088:13  */
  assign n6803_o = n6787_o ? 6'b000000 : n6792_o;
  /* control_fsm_rtl.vhd:2088:13  */
  assign n6806_o = n6787_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:2088:13  */
  assign n6808_o = n6787_o ? 4'b0000 : n6795_o;
  /* control_fsm_rtl.vhd:2088:13  */
  assign n6810_o = n6787_o ? 3'b000 : n6798_o;
  /* control_fsm_rtl.vhd:2088:13  */
  assign n6812_o = n6787_o ? 4'b0000 : n6801_o;
  /* control_fsm_rtl.vhd:2088:13  */
  assign n6815_o = n6787_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:2085:13  */
  assign n6817_o = n6785_o ? 6'b000000 : n6803_o;
  /* control_fsm_rtl.vhd:2085:13  */
  assign n6819_o = n6785_o ? 3'b010 : n6806_o;
  /* control_fsm_rtl.vhd:2085:13  */
  assign n6821_o = n6785_o ? 4'b0001 : n6808_o;
  /* control_fsm_rtl.vhd:2085:13  */
  assign n6823_o = n6785_o ? 3'b000 : n6810_o;
  /* control_fsm_rtl.vhd:2085:13  */
  assign n6825_o = n6785_o ? 4'b0000 : n6812_o;
  /* control_fsm_rtl.vhd:2085:13  */
  assign n6827_o = n6785_o ? 4'b0000 : n6815_o;
  /* control_fsm_rtl.vhd:2084:11  */
  assign n6829_o = s_instr_category == 7'b1101010;
  /* control_fsm_rtl.vhd:2101:21  */
  assign n6831_o = state == 3'b001;
  /* control_fsm_rtl.vhd:2104:24  */
  assign n6833_o = state == 3'b010;
  /* control_fsm_rtl.vhd:2104:13  */
  assign n6836_o = n6833_o ? 6'b101111 : 6'b000000;
  /* control_fsm_rtl.vhd:2104:13  */
  assign n6839_o = n6833_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:2104:13  */
  assign n6842_o = n6833_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:2104:13  */
  assign n6845_o = n6833_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:2101:13  */
  assign n6847_o = n6831_o ? 6'b000000 : n6836_o;
  /* control_fsm_rtl.vhd:2101:13  */
  assign n6850_o = n6831_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:2101:13  */
  assign n6852_o = n6831_o ? 4'b0000 : n6839_o;
  /* control_fsm_rtl.vhd:2101:13  */
  assign n6854_o = n6831_o ? 3'b000 : n6842_o;
  /* control_fsm_rtl.vhd:2101:13  */
  assign n6856_o = n6831_o ? 4'b0000 : n6845_o;
  /* control_fsm_rtl.vhd:2101:13  */
  assign n6859_o = n6831_o ? 4'b0111 : 4'b0000;
  /* control_fsm_rtl.vhd:2100:11  */
  assign n6861_o = s_instr_category == 7'b1101011;
  /* control_fsm_rtl.vhd:2114:21  */
  assign n6863_o = state == 3'b001;
  /* control_fsm_rtl.vhd:2117:24  */
  assign n6865_o = state == 3'b010;
  /* control_fsm_rtl.vhd:2117:13  */
  assign n6868_o = n6865_o ? 6'b110000 : 6'b000000;
  /* control_fsm_rtl.vhd:2117:13  */
  assign n6871_o = n6865_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:2117:13  */
  assign n6874_o = n6865_o ? 3'b010 : 3'b000;
  /* control_fsm_rtl.vhd:2117:13  */
  assign n6877_o = n6865_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:2114:13  */
  assign n6879_o = n6863_o ? 6'b000000 : n6868_o;
  /* control_fsm_rtl.vhd:2114:13  */
  assign n6882_o = n6863_o ? 3'b010 : 3'b001;
  /* control_fsm_rtl.vhd:2114:13  */
  assign n6884_o = n6863_o ? 4'b0001 : n6871_o;
  /* control_fsm_rtl.vhd:2114:13  */
  assign n6886_o = n6863_o ? 3'b000 : n6874_o;
  /* control_fsm_rtl.vhd:2114:13  */
  assign n6888_o = n6863_o ? 4'b0000 : n6877_o;
  /* control_fsm_rtl.vhd:2113:11  */
  assign n6890_o = s_instr_category == 7'b1101100;
  /* control_fsm_rtl.vhd:2127:21  */
  assign n6892_o = state == 3'b001;
  /* control_fsm_rtl.vhd:2130:24  */
  assign n6894_o = state == 3'b010;
  /* control_fsm_rtl.vhd:2133:24  */
  assign n6896_o = state == 3'b011;
  /* control_fsm_rtl.vhd:2133:13  */
  assign n6899_o = n6896_o ? 6'b101111 : 6'b000000;
  /* control_fsm_rtl.vhd:2133:13  */
  assign n6902_o = n6896_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:2133:13  */
  assign n6905_o = n6896_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:2133:13  */
  assign n6908_o = n6896_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:2133:13  */
  assign n6911_o = n6896_o ? 4'b1000 : 4'b0000;
  /* control_fsm_rtl.vhd:2130:13  */
  assign n6913_o = n6894_o ? 6'b000000 : n6899_o;
  /* control_fsm_rtl.vhd:2130:13  */
  assign n6916_o = n6894_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:2130:13  */
  assign n6918_o = n6894_o ? 4'b0000 : n6902_o;
  /* control_fsm_rtl.vhd:2130:13  */
  assign n6920_o = n6894_o ? 3'b000 : n6905_o;
  /* control_fsm_rtl.vhd:2130:13  */
  assign n6922_o = n6894_o ? 4'b0000 : n6908_o;
  /* control_fsm_rtl.vhd:2130:13  */
  assign n6924_o = n6894_o ? 4'b1000 : n6911_o;
  /* control_fsm_rtl.vhd:2127:13  */
  assign n6926_o = n6892_o ? 6'b000000 : n6913_o;
  /* control_fsm_rtl.vhd:2127:13  */
  assign n6928_o = n6892_o ? 3'b010 : n6916_o;
  /* control_fsm_rtl.vhd:2127:13  */
  assign n6930_o = n6892_o ? 4'b0001 : n6918_o;
  /* control_fsm_rtl.vhd:2127:13  */
  assign n6932_o = n6892_o ? 3'b000 : n6920_o;
  /* control_fsm_rtl.vhd:2127:13  */
  assign n6934_o = n6892_o ? 4'b0000 : n6922_o;
  /* control_fsm_rtl.vhd:2127:13  */
  assign n6936_o = n6892_o ? 4'b0000 : n6924_o;
  /* control_fsm_rtl.vhd:2126:11  */
  assign n6938_o = s_instr_category == 7'b1101101;
  /* control_fsm_rtl.vhd:2145:21  */
  assign n6940_o = state == 3'b001;
  /* control_fsm_rtl.vhd:2148:24  */
  assign n6942_o = state == 3'b010;
  /* control_fsm_rtl.vhd:2153:24  */
  assign n6944_o = state == 3'b011;
  /* control_fsm_rtl.vhd:2153:13  */
  assign n6947_o = n6944_o ? 6'b110001 : 6'b000000;
  /* control_fsm_rtl.vhd:2153:13  */
  assign n6950_o = n6944_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:2153:13  */
  assign n6953_o = n6944_o ? 3'b100 : 3'b000;
  /* control_fsm_rtl.vhd:2153:13  */
  assign n6956_o = n6944_o ? 4'b0011 : 4'b0000;
  /* control_fsm_rtl.vhd:2153:13  */
  assign n6959_o = n6944_o ? 4'b1010 : 4'b0000;
  /* control_fsm_rtl.vhd:2148:13  */
  assign n6961_o = n6942_o ? 6'b000000 : n6947_o;
  /* control_fsm_rtl.vhd:2148:13  */
  assign n6964_o = n6942_o ? 3'b011 : 3'b001;
  /* control_fsm_rtl.vhd:2148:13  */
  assign n6966_o = n6942_o ? 4'b0001 : n6950_o;
  /* control_fsm_rtl.vhd:2148:13  */
  assign n6968_o = n6942_o ? 3'b000 : n6953_o;
  /* control_fsm_rtl.vhd:2148:13  */
  assign n6970_o = n6942_o ? 4'b0000 : n6956_o;
  /* control_fsm_rtl.vhd:2148:13  */
  assign n6972_o = n6942_o ? 4'b1000 : n6959_o;
  /* control_fsm_rtl.vhd:2148:13  */
  assign n6975_o = n6942_o ? 4'b0001 : 4'b0000;
  /* control_fsm_rtl.vhd:2145:13  */
  assign n6977_o = n6940_o ? 6'b000000 : n6961_o;
  /* control_fsm_rtl.vhd:2145:13  */
  assign n6979_o = n6940_o ? 3'b010 : n6964_o;
  /* control_fsm_rtl.vhd:2145:13  */
  assign n6981_o = n6940_o ? 4'b0001 : n6966_o;
  /* control_fsm_rtl.vhd:2145:13  */
  assign n6983_o = n6940_o ? 3'b000 : n6968_o;
  /* control_fsm_rtl.vhd:2145:13  */
  assign n6985_o = n6940_o ? 4'b0000 : n6970_o;
  /* control_fsm_rtl.vhd:2145:13  */
  assign n6987_o = n6940_o ? 4'b0000 : n6972_o;
  /* control_fsm_rtl.vhd:2145:13  */
  assign n6989_o = n6940_o ? 4'b0000 : n6975_o;
  /* control_fsm_rtl.vhd:2144:11  */
  assign n6991_o = s_instr_category == 7'b1101110;
  assign n6992_o = {n6991_o, n6938_o, n6890_o, n6861_o, n6829_o, n6783_o, n6751_o, n6707_o, n6663_o, n6605_o, n6561_o, n6559_o, n6530_o, n6498_o, n6452_o, n6420_o, n6406_o, n6377_o, n6375_o, n6373_o, n6371_o, n6369_o, n6367_o, n6270_o, n6233_o, n6192_o, n6163_o, n6124_o, n6085_o, n6032_o, n5984_o, n5955_o, n5923_o, n5877_o, n5845_o, n5843_o, n5795_o, n5754_o, n5725_o, n5686_o, n5684_o, n5682_o, n5655_o, n5628_o, n5601_o, n5574_o, n5545_o, n5504_o, n5502_o, n5456_o, n5427_o, n5386_o, n5357_o, n5328_o, n5296_o, n5252_o, n5250_o, n5226_o, n5199_o, n5160_o, n5133_o, n5108_o, n5059_o, n5041_o, n5023_o, n5006_o, n4978_o, n4976_o, n4960_o, n4919_o, n4892_o, n4815_o, n4781_o, n4733_o, n4699_o, n4697_o, n4639_o, n4597_o, n4549_o, n4515_o, n4467_o, n4433_o, n4431_o, n4429_o, n4388_o, n4386_o, n4384_o, n4360_o, n4358_o, n4356_o, n4293_o, n4230_o, n4167_o, n4112_o, n4073_o, n4034_o, n3981_o, n3933_o, n3904_o, n3872_o, n3826_o, n3794_o, n3777_o, n3748_o, n3716_o, n3670_o, n3638_o, n3609_o, n3577_o, n3531_o, n3499_o};
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6977_o;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6926_o;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6879_o;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6847_o;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6817_o;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6769_o;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6548_o;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6516_o;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6486_o;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6438_o;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b110101;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b110100;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b110011;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b110010;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6071_o;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n6020_o;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n5973_o;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n5941_o;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n5911_o;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n5863_o;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = n5831_o;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7002_o = n4878_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7002_o = n4802_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7002_o = n4769_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7002_o = n4720_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7002_o = 6'b111110;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7002_o = n4683_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7002_o = n4623_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7002_o = n4585_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7002_o = n4536_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7002_o = n4503_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7002_o = n4454_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7002_o = 6'b111000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7002_o = 6'b100000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7002_o = 6'b110110;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7002_o = n4340_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7002_o = n4277_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7002_o = n4214_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7002_o = n4155_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7002_o = n4020_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7002_o = n3969_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7002_o = n3922_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7002_o = n3890_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7002_o = n3860_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7002_o = n3812_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7002_o = 6'b000000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7002_o = n3766_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7002_o = n3734_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7002_o = n3704_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7002_o = n3656_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7002_o = n3627_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7002_o = n3595_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7002_o = n3565_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7002_o = n3517_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7002_o = 6'b000000;
      default: n7002_o = 6'b000000;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6979_o;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6928_o;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6882_o;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6850_o;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6819_o;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6772_o;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6738_o;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6695_o;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6651_o;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6593_o;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6551_o;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6519_o;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6488_o;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6441_o;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6416_o;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6396_o;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6345_o;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6260_o;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6223_o;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6182_o;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6153_o;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6114_o;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6073_o;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n6022_o;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5976_o;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5944_o;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5913_o;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5866_o;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5833_o;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5785_o;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5744_o;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5715_o;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5671_o;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5644_o;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5617_o;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5590_o;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5564_o;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7023_o = n5535_o;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7023_o = n5490_o;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7023_o = n5446_o;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7023_o = n5417_o;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7023_o = n5376_o;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7023_o = n5347_o;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7023_o = n5315_o;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7023_o = n5283_o;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7023_o = n5242_o;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7023_o = n5215_o;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7023_o = n5189_o;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7023_o = n5149_o;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7023_o = n5127_o;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7023_o = n5093_o;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7023_o = n5055_o;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7023_o = n5037_o;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7023_o = n5019_o;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7023_o = n5000_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7023_o = n4972_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7023_o = n4950_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7023_o = n4913_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7023_o = n4880_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7023_o = n4805_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7023_o = n4771_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7023_o = n4723_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7023_o = n4685_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7023_o = n4626_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7023_o = n4587_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7023_o = n4539_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7023_o = n4505_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7023_o = n4457_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7023_o = n4419_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7023_o = n4376_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7023_o = 3'b001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7023_o = n4342_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7023_o = n4279_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7023_o = n4216_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7023_o = n4157_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7023_o = n4102_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7023_o = n4063_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7023_o = n4022_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7023_o = n3971_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7023_o = n3925_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7023_o = n3893_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7023_o = n3862_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7023_o = n3815_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7023_o = n3787_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7023_o = n3769_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7023_o = n3737_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7023_o = n3706_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7023_o = n3659_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7023_o = n3630_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7023_o = n3598_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7023_o = n3567_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7023_o = n3520_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7023_o = n3486_o;
      default: n7023_o = 3'b001;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6981_o;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6930_o;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6884_o;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6852_o;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6821_o;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6774_o;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6740_o;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6697_o;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6653_o;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6595_o;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6553_o;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6521_o;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6490_o;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6443_o;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6418_o;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6398_o;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6347_o;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6262_o;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6225_o;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6184_o;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6155_o;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6116_o;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6075_o;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n6024_o;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5978_o;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5946_o;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5915_o;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5868_o;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5835_o;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5787_o;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5746_o;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5717_o;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5673_o;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5646_o;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5619_o;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5592_o;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5566_o;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7044_o = n5537_o;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7044_o = n5492_o;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7044_o = n5448_o;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7044_o = n5419_o;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7044_o = n5378_o;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7044_o = n5349_o;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7044_o = n5317_o;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7044_o = n5285_o;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7044_o = n5244_o;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7044_o = n5217_o;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7044_o = n5191_o;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7044_o = n5151_o;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7044_o = n5129_o;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7044_o = n5095_o;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7044_o = n5057_o;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7044_o = n5039_o;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7044_o = n5021_o;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7044_o = n5002_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7044_o = 4'b0101;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7044_o = n4974_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7044_o = n4952_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7044_o = n4915_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7044_o = n4882_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7044_o = n4807_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7044_o = n4773_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7044_o = n4725_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7044_o = n4687_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7044_o = n4628_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7044_o = n4589_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7044_o = n4541_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7044_o = n4507_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7044_o = n4459_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7044_o = n4421_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7044_o = n4378_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7044_o = 4'b0001;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7044_o = n4344_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7044_o = n4281_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7044_o = n4218_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7044_o = n4159_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7044_o = n4104_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7044_o = n4065_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7044_o = n4024_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7044_o = n3973_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7044_o = n3927_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7044_o = n3895_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7044_o = n3864_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7044_o = n3817_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7044_o = n3789_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7044_o = n3771_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7044_o = n3739_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7044_o = n3708_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7044_o = n3661_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7044_o = n3632_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7044_o = n3600_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7044_o = n3569_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7044_o = n3522_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7044_o = n3488_o;
      default: n7044_o = 4'b0000;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6983_o;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6932_o;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6886_o;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6854_o;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6823_o;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6776_o;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6742_o;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6699_o;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6655_o;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6597_o;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = 3'b010;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6555_o;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6523_o;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6492_o;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6445_o;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6400_o;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = 3'b110;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = 3'b111;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = 3'b010;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = 3'b111;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = 3'b010;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6349_o;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6264_o;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6227_o;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6186_o;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6157_o;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6118_o;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6077_o;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n6026_o;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5980_o;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5948_o;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5917_o;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5870_o;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5837_o;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5789_o;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5748_o;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5719_o;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5675_o;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5648_o;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5621_o;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5594_o;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5568_o;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7061_o = n5539_o;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7061_o = 3'b100;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7061_o = n5494_o;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7061_o = n5450_o;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7061_o = n5421_o;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7061_o = n5380_o;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7061_o = n5351_o;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7061_o = n5319_o;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7061_o = n5287_o;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7061_o = 3'b100;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7061_o = n5246_o;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7061_o = n5219_o;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7061_o = n5193_o;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7061_o = n5153_o;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7061_o = n5097_o;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7061_o = n4954_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7061_o = n4884_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7061_o = n4809_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7061_o = n4775_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7061_o = n4727_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7061_o = 3'b010;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7061_o = n4689_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7061_o = n4630_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7061_o = n4591_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7061_o = n4543_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7061_o = n4509_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7061_o = n4461_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7061_o = 3'b010;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7061_o = 3'b111;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7061_o = n4423_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7061_o = 3'b110;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7061_o = 3'b010;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7061_o = n4380_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7061_o = 3'b110;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7061_o = 3'b010;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7061_o = n4346_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7061_o = n4283_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7061_o = n4220_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7061_o = n4161_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7061_o = n4106_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7061_o = n4067_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7061_o = n4026_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7061_o = n3975_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7061_o = n3929_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7061_o = n3897_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7061_o = n3866_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7061_o = n3819_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7061_o = 3'b000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7061_o = n3773_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7061_o = n3741_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7061_o = n3710_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7061_o = n3663_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7061_o = n3634_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7061_o = n3602_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7061_o = n3571_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7061_o = n3524_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7061_o = n3490_o;
      default: n7061_o = 3'b000;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6985_o;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6934_o;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6888_o;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6856_o;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6825_o;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6778_o;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6744_o;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6701_o;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6657_o;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6599_o;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0111;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6557_o;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6525_o;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6494_o;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6447_o;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0011;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0011;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0011;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0011;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6229_o;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6188_o;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6079_o;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n6028_o;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5982_o;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5950_o;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5919_o;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5872_o;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5839_o;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5791_o;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5677_o;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5650_o;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5623_o;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5596_o;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5570_o;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7075_o = n5541_o;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0110;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7075_o = n5496_o;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7075_o = n5452_o;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7075_o = n5423_o;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7075_o = n5382_o;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7075_o = n5353_o;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7075_o = n5321_o;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7075_o = n5289_o;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7075_o = 4'b0110;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7075_o = n5248_o;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7075_o = n5221_o;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7075_o = n5195_o;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7075_o = n5155_o;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7075_o = n5099_o;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7075_o = n4886_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7075_o = n4811_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7075_o = n4777_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7075_o = n4729_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7075_o = 4'b0011;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7075_o = n4691_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7075_o = n4632_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7075_o = n4593_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7075_o = n4545_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7075_o = n4511_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7075_o = n4463_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7075_o = 4'b0011;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7075_o = 4'b0011;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7075_o = 4'b0011;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7075_o = n4028_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7075_o = n3977_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7075_o = n3931_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7075_o = n3899_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7075_o = n3868_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7075_o = n3821_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7075_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7075_o = n3775_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7075_o = n3743_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7075_o = n3712_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7075_o = n3665_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7075_o = n3636_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7075_o = n3604_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7075_o = n3573_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7075_o = n3526_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7075_o = n3492_o;
      default: n7075_o = 4'b0000;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = n6402_o;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b1011;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = n6159_o;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = n6120_o;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = n5750_o;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = n5721_o;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7080_o = n4425_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7080_o = 4'b0101;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7080_o = n4348_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7080_o = n4285_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7080_o = n4222_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7080_o = n4163_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7080_o = n4108_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7080_o = n4069_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7080_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7080_o = 4'b0000;
      default: n7080_o = 4'b0000;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6987_o;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6936_o;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6859_o;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6827_o;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6781_o;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6746_o;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6703_o;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6659_o;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6601_o;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6528_o;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6496_o;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6450_o;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6404_o;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b1011;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6351_o;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6266_o;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6231_o;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6190_o;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6161_o;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6122_o;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6081_o;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n6030_o;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n5953_o;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n5921_o;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n5875_o;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n5841_o;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n5793_o;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n5752_o;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = n5723_o;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7087_o = n5572_o;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7087_o = n5543_o;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0111;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7087_o = n5498_o;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7087_o = n5454_o;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7087_o = n5425_o;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7087_o = n5384_o;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7087_o = n5355_o;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7087_o = n5323_o;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7087_o = n5291_o;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0110;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7087_o = n5224_o;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7087_o = n5197_o;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7087_o = n5158_o;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7087_o = n5101_o;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7087_o = n5004_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7087_o = n4956_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7087_o = n4917_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7087_o = n4888_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7087_o = n4813_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7087_o = n4779_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7087_o = n4731_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7087_o = n4693_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7087_o = n4634_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7087_o = n4595_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7087_o = n4547_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7087_o = n4513_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7087_o = n4465_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7087_o = n4427_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7087_o = 4'b1011;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7087_o = n4382_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7087_o = 4'b1011;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7087_o = n4350_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7087_o = n4287_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7087_o = n4224_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7087_o = n4165_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7087_o = n4110_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7087_o = n4071_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7087_o = n4030_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7087_o = n3979_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7087_o = n3902_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7087_o = n3870_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7087_o = n3824_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7087_o = n3746_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7087_o = n3714_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7087_o = n3668_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7087_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7087_o = n3607_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7087_o = n3575_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7087_o = n3529_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7087_o = n3494_o;
      default: n7087_o = 4'b0000;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b01;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b10;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7091_o = n5680_o;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7091_o = n5653_o;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7091_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7091_o = 2'b00;
      default: n7091_o = 2'b00;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b1;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b1;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7095_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7095_o = 1'b0;
      default: n7095_o = 1'b0;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = n6989_o;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = n6749_o;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = n6705_o;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = n6661_o;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = n6603_o;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = n6353_o;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = n6268_o;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = n6083_o;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7097_o = n5500_o;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7097_o = n5326_o;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7097_o = n5294_o;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7097_o = n5131_o;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7097_o = n5103_o;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7097_o = n4958_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7097_o = n4890_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7097_o = n4695_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7097_o = n4637_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7097_o = n4352_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7097_o = n4289_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7097_o = n4226_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7097_o = n4032_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7097_o = 4'b0000;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7097_o = 4'b0000;
      default: n7097_o = 4'b0000;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7099_o = n5626_o;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7099_o = n5599_o;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7099_o = n5106_o;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7099_o = n3792_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7099_o = 2'b00;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7099_o = n3497_o;
      default: n7099_o = 2'b00;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7101_o = n4354_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7101_o = n4291_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7101_o = n4228_o;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7101_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7101_o = 1'b0;
      default: n7101_o = 1'b0;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = n6355_o;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7103_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7103_o = 1'b0;
      default: n7103_o = 1'b0;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = n6357_o;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7105_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7105_o = 1'b0;
      default: n7105_o = 1'b0;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = n6359_o;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7107_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7107_o = 1'b0;
      default: n7107_o = 1'b0;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = n6361_o;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7109_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7109_o = 1'b0;
      default: n7109_o = 1'b0;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = n6363_o;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7111_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7111_o = 1'b0;
      default: n7111_o = 1'b0;
    endcase
  /* control_fsm_rtl.vhd:439:9  */
  always @*
    case (n6992_o)
      111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = n6365_o;
      111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7113_o = 1'b0;
      111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7113_o = 1'b0;
      default: n7113_o = 1'b0;
    endcase
  /* control_fsm_rtl.vhd:340:7  */
  assign n7115_o = n3134_o ? 6'b000000 : n7002_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7116_o = n3134_o ? n3428_o : n7023_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7117_o = n3134_o ? n3430_o : n7044_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7118_o = n3134_o ? n3432_o : n7061_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7119_o = n3134_o ? n3434_o : n7075_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7121_o = n3134_o ? 4'b0000 : n7080_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7122_o = n3134_o ? n3436_o : n7087_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7124_o = n3134_o ? 2'b00 : n7091_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7126_o = n3134_o ? 1'b0 : n7095_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7127_o = n3134_o ? n3438_o : n7097_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7129_o = n3134_o ? 2'b00 : n7099_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7131_o = n3134_o ? 1'b0 : n7101_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7133_o = n3134_o ? n3441_o : 1'b0;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7135_o = n3134_o ? n3443_o : 1'b0;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7137_o = n3134_o ? n3445_o : 1'b0;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7138_o = n3134_o ? n3447_o : n7103_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7140_o = n3134_o ? n3449_o : 1'b0;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7141_o = n3134_o ? n3451_o : n7105_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7143_o = n3134_o ? n3453_o : 1'b0;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7145_o = n3134_o ? n3455_o : 1'b0;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7147_o = n3134_o ? n3457_o : 1'b0;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7149_o = n3134_o ? n3459_o : 1'b0;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7150_o = n3134_o ? n3461_o : n7107_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7151_o = n3134_o ? n3463_o : n7109_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7152_o = n3134_o ? n3465_o : n7111_o;
  /* control_fsm_rtl.vhd:340:7  */
  assign n7153_o = n3134_o ? n3467_o : n7113_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7155_o = n3125_o ? 6'b000000 : n7115_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7158_o = n3125_o ? 3'b001 : n7116_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7161_o = n3125_o ? 4'b0000 : n7117_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7164_o = n3125_o ? 3'b000 : n7118_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7167_o = n3125_o ? 4'b0000 : n7119_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7170_o = n3125_o ? 4'b0000 : n7121_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7173_o = n3125_o ? 4'b0000 : n7122_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7176_o = n3125_o ? 2'b00 : n7124_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7179_o = n3125_o ? 1'b0 : n7126_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7182_o = n3125_o ? 4'b0000 : n7127_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7185_o = n3125_o ? 2'b00 : n7129_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7188_o = n3125_o ? 1'b0 : n7131_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7191_o = n3125_o ? 1'b0 : n7133_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7194_o = n3125_o ? 1'b0 : n7135_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7197_o = n3125_o ? 1'b0 : n7137_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7200_o = n3125_o ? 1'b0 : n7138_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7203_o = n3125_o ? 1'b0 : n7140_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7206_o = n3125_o ? 1'b0 : n7141_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7209_o = n3125_o ? 1'b0 : n7143_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7212_o = n3125_o ? 1'b0 : n7145_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7215_o = n3125_o ? 1'b0 : n7147_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7218_o = n3125_o ? 1'b0 : n7149_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7221_o = n3125_o ? 1'b0 : n7150_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7224_o = n3125_o ? 1'b0 : n7151_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7227_o = n3125_o ? 1'b0 : n7152_o;
  /* control_fsm_rtl.vhd:334:5  */
  assign n7230_o = n3125_o ? 1'b0 : n7153_o;
endmodule

module mc8051_tmrctr
  (input  clk,
   input  cen,
   input  reset,
   input  int0_i,
   input  int1_i,
   input  t0_i,
   input  t1_i,
   input  [7:0] tmod_i,
   input  tcon_tr0_i,
   input  tcon_tr1_i,
   input  [7:0] reload_i,
   input  wt_en_i,
   input  [1:0] wt_i,
   output [7:0] th0_o,
   output [7:0] tl0_o,
   output [7:0] th1_o,
   output [7:0] tl1_o,
   output tf0_o,
   output tf1_o);
  wire [3:0] s_pre_count;
  wire s_count_enable;
  wire [15:0] s_count0;
  wire [7:0] s_countl0;
  wire [7:0] s_counth0;
  wire [15:0] s_count1;
  wire [7:0] s_countl1;
  wire [7:0] s_counth1;
  wire s_gate0;
  wire s_gate1;
  wire s_c_t0;
  wire s_c_t1;
  wire s_tmr_ctr0_en;
  wire s_tmr_ctr1_en;
  wire [1:0] s_mode0;
  wire [1:0] s_mode1;
  wire s_tf0;
  wire s_tf1;
  wire s_t0ff0;
  wire s_t0ff1;
  wire s_t0ff2;
  wire s_t1ff0;
  wire s_t1ff1;
  wire s_t1ff2;
  wire s_ext_edge0;
  wire s_ext_edge1;
  wire [1:0] s_int0_sync;
  wire [1:0] s_int1_sync;
  wire n1970_o;
  wire n1971_o;
  wire n1972_o;
  wire n1973_o;
  wire n1974_o;
  wire n1975_o;
  wire n1976_o;
  wire n1977_o;
  wire n1978_o;
  wire n1979_o;
  wire n1980_o;
  wire n1981_o;
  wire n1982_o;
  wire n1983_o;
  wire n1984_o;
  wire n1986_o;
  wire n1987_o;
  wire n1988_o;
  wire n1989_o;
  wire n1990_o;
  wire n1991_o;
  wire [7:0] n1992_o;
  wire [7:0] n1993_o;
  wire [7:0] n1994_o;
  wire [7:0] n1995_o;
  wire n1998_o;
  wire n1999_o;
  wire [3:0] n2006_o;
  wire n2008_o;
  wire [3:0] n2010_o;
  wire n2011_o;
  wire n2012_o;
  wire [1:0] n2014_o;
  wire [1:0] n2016_o;
  wire n2026_o;
  wire n2027_o;
  wire n2028_o;
  wire n2032_o;
  wire n2035_o;
  wire n2039_o;
  wire n2040_o;
  wire n2041_o;
  wire n2053_o;
  wire n2054_o;
  wire n2055_o;
  wire n2059_o;
  wire n2062_o;
  wire n2066_o;
  wire n2067_o;
  wire n2068_o;
  wire n2082_o;
  wire n2083_o;
  wire n2084_o;
  wire n2086_o;
  wire n2089_o;
  wire n2091_o;
  wire n2093_o;
  wire n2095_o;
  wire n2097_o;
  wire n2098_o;
  wire n2099_o;
  wire n2101_o;
  wire [7:0] n2104_o;
  wire [7:0] n2106_o;
  wire n2108_o;
  wire [7:0] n2111_o;
  wire [7:0] n2113_o;
  wire [7:0] n2114_o;
  wire [7:0] n2115_o;
  wire [7:0] n2116_o;
  wire n2117_o;
  wire [7:0] n2118_o;
  wire n2120_o;
  wire n2121_o;
  wire n2122_o;
  wire n2124_o;
  wire n2126_o;
  wire [7:0] n2129_o;
  wire [7:0] n2130_o;
  wire [7:0] n2132_o;
  wire n2134_o;
  wire n2136_o;
  wire [7:0] n2139_o;
  wire [7:0] n2140_o;
  wire [7:0] n2142_o;
  wire [7:0] n2143_o;
  wire [7:0] n2144_o;
  wire [7:0] n2145_o;
  wire n2146_o;
  wire [7:0] n2147_o;
  wire n2149_o;
  wire n2150_o;
  wire n2151_o;
  wire n2152_o;
  wire n2154_o;
  wire n2157_o;
  wire n2159_o;
  wire n2161_o;
  wire n2163_o;
  wire n2165_o;
  wire n2166_o;
  wire n2167_o;
  wire n2169_o;
  wire [7:0] n2172_o;
  wire [7:0] n2174_o;
  wire n2176_o;
  wire [7:0] n2179_o;
  wire [7:0] n2181_o;
  wire [7:0] n2182_o;
  wire [7:0] n2183_o;
  wire [7:0] n2184_o;
  wire n2185_o;
  wire [7:0] n2186_o;
  wire n2188_o;
  wire n2189_o;
  wire n2190_o;
  wire n2192_o;
  wire n2194_o;
  wire [7:0] n2197_o;
  wire [7:0] n2198_o;
  wire [7:0] n2200_o;
  wire n2202_o;
  wire n2204_o;
  wire [7:0] n2207_o;
  wire [7:0] n2208_o;
  wire [7:0] n2210_o;
  wire [7:0] n2211_o;
  wire [7:0] n2212_o;
  wire [7:0] n2213_o;
  wire n2214_o;
  wire [7:0] n2215_o;
  wire n2217_o;
  wire n2218_o;
  wire n2219_o;
  wire n2220_o;
  wire [7:0] n2221_o;
  wire [15:0] n2222_o;
  wire n2224_o;
  wire n2227_o;
  wire n2229_o;
  wire n2231_o;
  wire n2233_o;
  wire n2235_o;
  wire n2236_o;
  wire n2237_o;
  wire n2239_o;
  wire [7:0] n2242_o;
  wire [7:0] n2243_o;
  wire n2245_o;
  wire [7:0] n2248_o;
  wire [7:0] n2249_o;
  wire [7:0] n2250_o;
  wire [7:0] n2251_o;
  wire [7:0] n2252_o;
  wire n2253_o;
  wire [7:0] n2254_o;
  wire n2256_o;
  wire n2257_o;
  wire [7:0] n2258_o;
  wire n2260_o;
  wire n2261_o;
  wire n2262_o;
  wire n2263_o;
  wire [7:0] n2264_o;
  wire [15:0] n2265_o;
  wire n2267_o;
  wire n2270_o;
  wire n2272_o;
  wire n2274_o;
  wire n2276_o;
  wire n2278_o;
  wire n2279_o;
  wire n2280_o;
  wire n2282_o;
  wire [7:0] n2285_o;
  wire [7:0] n2287_o;
  wire n2289_o;
  wire [7:0] n2292_o;
  wire [7:0] n2294_o;
  wire [7:0] n2295_o;
  wire [7:0] n2296_o;
  wire [7:0] n2297_o;
  wire n2298_o;
  wire [7:0] n2299_o;
  wire [7:0] n2300_o;
  wire n2302_o;
  wire n2305_o;
  wire n2307_o;
  wire n2309_o;
  wire n2311_o;
  wire n2312_o;
  wire n2314_o;
  wire [7:0] n2317_o;
  wire [7:0] n2319_o;
  wire [7:0] n2320_o;
  wire n2321_o;
  wire [7:0] n2322_o;
  wire n2324_o;
  wire [3:0] n2325_o;
  reg [7:0] n2326_o;
  reg [7:0] n2327_o;
  reg n2329_o;
  reg n2332_o;
  wire n2335_o;
  wire n2337_o;
  wire n2338_o;
  wire n2340_o;
  wire n2341_o;
  wire n2342_o;
  wire n2343_o;
  wire n2344_o;
  wire n2346_o;
  wire n2349_o;
  wire n2350_o;
  wire n2351_o;
  wire n2352_o;
  wire n2353_o;
  wire n2355_o;
  wire n2356_o;
  wire n2357_o;
  wire n2359_o;
  wire [7:0] n2362_o;
  wire [7:0] n2364_o;
  wire n2366_o;
  wire [7:0] n2369_o;
  wire [7:0] n2371_o;
  wire [7:0] n2372_o;
  wire [7:0] n2373_o;
  wire [7:0] n2374_o;
  wire n2375_o;
  wire [7:0] n2376_o;
  wire n2378_o;
  wire n2379_o;
  wire n2380_o;
  wire n2382_o;
  wire n2384_o;
  wire [7:0] n2387_o;
  wire [7:0] n2388_o;
  wire [7:0] n2390_o;
  wire n2392_o;
  wire n2394_o;
  wire [7:0] n2397_o;
  wire [7:0] n2398_o;
  wire [7:0] n2400_o;
  wire [7:0] n2401_o;
  wire [7:0] n2402_o;
  wire [7:0] n2403_o;
  wire n2404_o;
  wire [7:0] n2405_o;
  wire n2407_o;
  wire n2409_o;
  wire n2411_o;
  wire n2412_o;
  wire n2414_o;
  wire n2415_o;
  wire n2416_o;
  wire n2417_o;
  wire n2418_o;
  wire n2420_o;
  wire n2423_o;
  wire n2424_o;
  wire n2425_o;
  wire n2426_o;
  wire n2427_o;
  wire n2429_o;
  wire n2430_o;
  wire n2431_o;
  wire n2433_o;
  wire [7:0] n2436_o;
  wire [7:0] n2438_o;
  wire n2440_o;
  wire [7:0] n2443_o;
  wire [7:0] n2445_o;
  wire [7:0] n2446_o;
  wire [7:0] n2447_o;
  wire [7:0] n2448_o;
  wire n2449_o;
  wire [7:0] n2450_o;
  wire n2452_o;
  wire n2453_o;
  wire n2454_o;
  wire n2456_o;
  wire n2458_o;
  wire [7:0] n2461_o;
  wire [7:0] n2462_o;
  wire [7:0] n2464_o;
  wire n2466_o;
  wire n2468_o;
  wire [7:0] n2471_o;
  wire [7:0] n2472_o;
  wire [7:0] n2474_o;
  wire [7:0] n2475_o;
  wire [7:0] n2476_o;
  wire [7:0] n2477_o;
  wire n2478_o;
  wire [7:0] n2479_o;
  wire n2481_o;
  wire n2483_o;
  wire n2485_o;
  wire n2486_o;
  wire n2488_o;
  wire n2489_o;
  wire n2490_o;
  wire n2491_o;
  wire n2492_o;
  wire [7:0] n2493_o;
  wire [15:0] n2494_o;
  wire n2496_o;
  wire n2499_o;
  wire n2500_o;
  wire n2501_o;
  wire n2502_o;
  wire n2503_o;
  wire n2505_o;
  wire n2506_o;
  wire n2507_o;
  wire n2509_o;
  wire [7:0] n2512_o;
  wire [7:0] n2513_o;
  wire n2515_o;
  wire [7:0] n2518_o;
  wire [7:0] n2519_o;
  wire [7:0] n2520_o;
  wire [7:0] n2521_o;
  wire [7:0] n2522_o;
  wire n2523_o;
  wire [7:0] n2524_o;
  wire n2526_o;
  wire n2527_o;
  wire [7:0] n2528_o;
  wire n2530_o;
  wire n2532_o;
  wire n2533_o;
  wire [7:0] n2534_o;
  wire n2536_o;
  wire n2537_o;
  wire [7:0] n2538_o;
  wire n2540_o;
  wire [3:0] n2541_o;
  reg [7:0] n2542_o;
  reg [7:0] n2543_o;
  reg n2544_o;
  wire [3:0] n2564_o;
  reg [3:0] n2565_q;
  wire [15:0] n2566_o;
  wire [7:0] n2567_o;
  reg [7:0] n2568_q;
  wire [7:0] n2569_o;
  reg [7:0] n2570_q;
  wire [15:0] n2571_o;
  wire [7:0] n2572_o;
  reg [7:0] n2573_q;
  wire [7:0] n2574_o;
  reg [7:0] n2575_q;
  wire [1:0] n2576_o;
  wire [1:0] n2577_o;
  wire n2578_o;
  reg n2579_q;
  wire n2580_o;
  reg n2581_q;
  wire n2582_o;
  wire n2583_o;
  reg n2584_q;
  wire n2585_o;
  wire n2586_o;
  reg n2587_q;
  wire n2588_o;
  reg n2589_q;
  wire n2590_o;
  wire n2591_o;
  reg n2592_q;
  wire n2593_o;
  wire n2594_o;
  reg n2595_q;
  wire n2596_o;
  reg n2597_q;
  wire [1:0] n2598_o;
  reg [1:0] n2599_q;
  wire [1:0] n2600_o;
  reg [1:0] n2601_q;
  assign th0_o = n1992_o;
  assign tl0_o = n1993_o;
  assign th1_o = n1994_o;
  assign tl1_o = n1995_o;
  assign tf0_o = s_tf0;
  assign tf1_o = s_tf1;
  /* mc8051_tmrctr_rtl.vhd:67:10  */
  assign s_pre_count = n2565_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:68:10  */
  assign s_count_enable = n1999_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:72:10  */
  assign s_count0 = n2566_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:73:10  */
  assign s_countl0 = n2568_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:74:10  */
  assign s_counth0 = n2570_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:75:10  */
  assign s_count1 = n2571_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:76:10  */
  assign s_countl1 = n2573_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:77:10  */
  assign s_counth1 = n2575_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:78:10  */
  assign s_gate0 = n1970_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:79:10  */
  assign s_gate1 = n1974_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:80:10  */
  assign s_c_t0 = n1971_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:81:10  */
  assign s_c_t1 = n1975_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:82:10  */
  assign s_tmr_ctr0_en = n1981_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:83:10  */
  assign s_tmr_ctr1_en = n1987_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:84:10  */
  assign s_mode0 = n2576_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:85:10  */
  assign s_mode1 = n2577_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:86:10  */
  assign s_tf0 = n2579_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:87:10  */
  assign s_tf1 = n2581_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:88:10  */
  assign s_t0ff0 = n2584_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:89:10  */
  assign s_t0ff1 = n2587_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:90:10  */
  assign s_t0ff2 = n2589_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:91:10  */
  assign s_t1ff0 = n2592_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:92:10  */
  assign s_t1ff1 = n2595_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:93:10  */
  assign s_t1ff2 = n2597_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:94:10  */
  assign s_ext_edge0 = n2028_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:95:10  */
  assign s_ext_edge1 = n2055_o; // (signal)
  /* mc8051_tmrctr_rtl.vhd:96:10  */
  assign s_int0_sync = n2599_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:97:10  */
  assign s_int1_sync = n2601_q; // (signal)
  /* mc8051_tmrctr_rtl.vhd:103:20  */
  assign n1970_o = tmod_i[3];
  /* mc8051_tmrctr_rtl.vhd:104:20  */
  assign n1971_o = tmod_i[2];
  /* mc8051_tmrctr_rtl.vhd:105:23  */
  assign n1972_o = tmod_i[1];
  /* mc8051_tmrctr_rtl.vhd:106:23  */
  assign n1973_o = tmod_i[0];
  /* mc8051_tmrctr_rtl.vhd:108:20  */
  assign n1974_o = tmod_i[7];
  /* mc8051_tmrctr_rtl.vhd:109:20  */
  assign n1975_o = tmod_i[6];
  /* mc8051_tmrctr_rtl.vhd:110:23  */
  assign n1976_o = tmod_i[5];
  /* mc8051_tmrctr_rtl.vhd:111:23  */
  assign n1977_o = tmod_i[4];
  /* mc8051_tmrctr_rtl.vhd:114:36  */
  assign n1978_o = ~s_gate0;
  /* mc8051_tmrctr_rtl.vhd:114:63  */
  assign n1979_o = s_int0_sync[1];
  /* mc8051_tmrctr_rtl.vhd:114:49  */
  assign n1980_o = n1978_o | n1979_o;
  /* mc8051_tmrctr_rtl.vhd:114:31  */
  assign n1981_o = tcon_tr0_i & n1980_o;
  /* mc8051_tmrctr_rtl.vhd:115:21  */
  assign n1982_o = ~s_gate1;
  /* mc8051_tmrctr_rtl.vhd:115:48  */
  assign n1983_o = s_int1_sync[1];
  /* mc8051_tmrctr_rtl.vhd:115:34  */
  assign n1984_o = n1982_o | n1983_o;
  /* mc8051_tmrctr_rtl.vhd:116:55  */
  assign n1986_o = s_mode0 == 2'b11;
  /* mc8051_tmrctr_rtl.vhd:115:53  */
  assign n1987_o = n1986_o ? n1984_o : n1991_o;
  /* mc8051_tmrctr_rtl.vhd:117:36  */
  assign n1988_o = ~s_gate1;
  /* mc8051_tmrctr_rtl.vhd:117:63  */
  assign n1989_o = s_int1_sync[1];
  /* mc8051_tmrctr_rtl.vhd:117:49  */
  assign n1990_o = n1988_o | n1989_o;
  /* mc8051_tmrctr_rtl.vhd:117:31  */
  assign n1991_o = tcon_tr1_i & n1990_o;
  /* mc8051_tmrctr_rtl.vhd:124:37  */
  assign n1992_o = s_count0[15:8];
  /* mc8051_tmrctr_rtl.vhd:125:37  */
  assign n1993_o = s_count0[7:0];
  /* mc8051_tmrctr_rtl.vhd:126:37  */
  assign n1994_o = s_count1[15:8];
  /* mc8051_tmrctr_rtl.vhd:127:37  */
  assign n1995_o = s_count1[7:0];
  /* mc8051_tmrctr_rtl.vhd:135:42  */
  assign n1998_o = s_pre_count == 4'b1011;
  /* mc8051_tmrctr_rtl.vhd:135:25  */
  assign n1999_o = n1998_o ? 1'b1 : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:147:38  */
  assign n2006_o = s_pre_count + 4'b0001;
  /* mc8051_tmrctr_rtl.vhd:148:26  */
  assign n2008_o = s_pre_count == 4'b1011;
  /* mc8051_tmrctr_rtl.vhd:148:11  */
  assign n2010_o = n2008_o ? 4'b0000 : n2006_o;
  /* mc8051_tmrctr_rtl.vhd:152:40  */
  assign n2011_o = s_int0_sync[0];
  /* mc8051_tmrctr_rtl.vhd:154:40  */
  assign n2012_o = s_int1_sync[0];
  assign n2014_o = {n2011_o, int0_i};
  assign n2016_o = {n2012_o, int1_i};
  /* mc8051_tmrctr_rtl.vhd:166:36  */
  assign n2026_o = ~s_t0ff1;
  /* mc8051_tmrctr_rtl.vhd:166:42  */
  assign n2027_o = n2026_o & s_t0ff2;
  /* mc8051_tmrctr_rtl.vhd:166:22  */
  assign n2028_o = n2027_o ? 1'b1 : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:178:36  */
  assign n2032_o = cen & n2041_o;
  /* mc8051_tmrctr_rtl.vhd:179:26  */
  assign n2035_o = s_pre_count == 4'b0110;
  /* mc8051_tmrctr_rtl.vhd:179:11  */
  assign n2039_o = n2035_o & s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:179:11  */
  assign n2040_o = n2035_o & s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:179:11  */
  assign n2041_o = n2035_o & s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:191:36  */
  assign n2053_o = ~s_t1ff1;
  /* mc8051_tmrctr_rtl.vhd:191:42  */
  assign n2054_o = n2053_o & s_t1ff2;
  /* mc8051_tmrctr_rtl.vhd:191:22  */
  assign n2055_o = n2054_o ? 1'b1 : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:202:36  */
  assign n2059_o = cen & n2068_o;
  /* mc8051_tmrctr_rtl.vhd:203:26  */
  assign n2062_o = s_pre_count == 4'b0110;
  /* mc8051_tmrctr_rtl.vhd:203:11  */
  assign n2066_o = n2062_o & s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:203:11  */
  assign n2067_o = n2062_o & s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:203:11  */
  assign n2068_o = n2062_o & s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:254:23  */
  assign n2082_o = ~s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:254:51  */
  assign n2083_o = s_ext_edge0 & s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:254:29  */
  assign n2084_o = n2082_o | n2083_o;
  /* mc8051_tmrctr_rtl.vhd:255:27  */
  assign n2086_o = s_count0 == 16'b1111111100011111;
  /* mc8051_tmrctr_rtl.vhd:255:15  */
  assign n2089_o = n2086_o ? 1'b1 : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:254:13  */
  assign n2091_o = n2084_o ? n2089_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:253:11  */
  assign n2093_o = s_count_enable ? n2091_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:252:9  */
  assign n2095_o = s_tmr_ctr0_en ? n2093_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:265:17  */
  assign n2097_o = wt_i == 2'b00;
  /* mc8051_tmrctr_rtl.vhd:265:24  */
  assign n2098_o = n2097_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:270:25  */
  assign n2099_o = ~s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:271:30  */
  assign n2101_o = s_countl0 == 8'b00011111;
  /* mc8051_tmrctr_rtl.vhd:274:42  */
  assign n2104_o = s_countl0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:271:17  */
  assign n2106_o = n2101_o ? 8'b00000000 : n2104_o;
  /* mc8051_tmrctr_rtl.vhd:278:32  */
  assign n2108_o = s_countl0 == 8'b00011111;
  /* mc8051_tmrctr_rtl.vhd:281:44  */
  assign n2111_o = s_countl0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:278:19  */
  assign n2113_o = n2108_o ? 8'b00000000 : n2111_o;
  /* mc8051_tmrctr_rtl.vhd:277:17  */
  assign n2114_o = s_ext_edge0 ? n2113_o : s_countl0;
  /* mc8051_tmrctr_rtl.vhd:270:15  */
  assign n2115_o = n2099_o ? n2106_o : n2114_o;
  /* mc8051_tmrctr_rtl.vhd:268:11  */
  assign n2116_o = n2117_o ? n2115_o : s_countl0;
  /* mc8051_tmrctr_rtl.vhd:268:11  */
  assign n2117_o = s_tmr_ctr0_en & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:265:9  */
  assign n2118_o = n2098_o ? reload_i : n2116_o;
  /* mc8051_tmrctr_rtl.vhd:290:17  */
  assign n2120_o = wt_i == 2'b10;
  /* mc8051_tmrctr_rtl.vhd:290:24  */
  assign n2121_o = n2120_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:295:25  */
  assign n2122_o = ~s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:296:29  */
  assign n2124_o = s_count0 == 16'b1111111100011111;
  /* mc8051_tmrctr_rtl.vhd:299:32  */
  assign n2126_o = s_countl0 == 8'b00011111;
  /* mc8051_tmrctr_rtl.vhd:300:44  */
  assign n2129_o = s_counth0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:299:19  */
  assign n2130_o = n2126_o ? n2129_o : s_counth0;
  /* mc8051_tmrctr_rtl.vhd:296:17  */
  assign n2132_o = n2124_o ? 8'b00000000 : n2130_o;
  /* mc8051_tmrctr_rtl.vhd:305:31  */
  assign n2134_o = s_count0 == 16'b1111111100011111;
  /* mc8051_tmrctr_rtl.vhd:308:34  */
  assign n2136_o = s_countl0 == 8'b00011111;
  /* mc8051_tmrctr_rtl.vhd:309:46  */
  assign n2139_o = s_counth0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:308:21  */
  assign n2140_o = n2136_o ? n2139_o : s_counth0;
  /* mc8051_tmrctr_rtl.vhd:305:19  */
  assign n2142_o = n2134_o ? 8'b00000000 : n2140_o;
  /* mc8051_tmrctr_rtl.vhd:304:17  */
  assign n2143_o = s_ext_edge0 ? n2142_o : s_counth0;
  /* mc8051_tmrctr_rtl.vhd:295:15  */
  assign n2144_o = n2122_o ? n2132_o : n2143_o;
  /* mc8051_tmrctr_rtl.vhd:293:11  */
  assign n2145_o = n2146_o ? n2144_o : s_counth0;
  /* mc8051_tmrctr_rtl.vhd:293:11  */
  assign n2146_o = s_tmr_ctr0_en & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:290:9  */
  assign n2147_o = n2121_o ? reload_i : n2145_o;
  /* mc8051_tmrctr_rtl.vhd:249:9  */
  assign n2149_o = s_mode0 == 2'b00;
  /* mc8051_tmrctr_rtl.vhd:326:23  */
  assign n2150_o = ~s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:326:51  */
  assign n2151_o = s_ext_edge0 & s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:326:29  */
  assign n2152_o = n2150_o | n2151_o;
  /* mc8051_tmrctr_rtl.vhd:327:27  */
  assign n2154_o = s_count0 == 16'b1111111111111111;
  /* mc8051_tmrctr_rtl.vhd:327:15  */
  assign n2157_o = n2154_o ? 1'b1 : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:326:13  */
  assign n2159_o = n2152_o ? n2157_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:325:11  */
  assign n2161_o = s_count_enable ? n2159_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:324:9  */
  assign n2163_o = s_tmr_ctr0_en ? n2161_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:337:17  */
  assign n2165_o = wt_i == 2'b00;
  /* mc8051_tmrctr_rtl.vhd:337:24  */
  assign n2166_o = n2165_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:342:25  */
  assign n2167_o = ~s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:343:29  */
  assign n2169_o = s_count0 == 16'b1111111111111111;
  /* mc8051_tmrctr_rtl.vhd:346:42  */
  assign n2172_o = s_countl0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:343:17  */
  assign n2174_o = n2169_o ? 8'b00000000 : n2172_o;
  /* mc8051_tmrctr_rtl.vhd:350:31  */
  assign n2176_o = s_count0 == 16'b1111111111111111;
  /* mc8051_tmrctr_rtl.vhd:353:44  */
  assign n2179_o = s_countl0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:350:19  */
  assign n2181_o = n2176_o ? 8'b00000000 : n2179_o;
  /* mc8051_tmrctr_rtl.vhd:349:17  */
  assign n2182_o = s_ext_edge0 ? n2181_o : s_countl0;
  /* mc8051_tmrctr_rtl.vhd:342:15  */
  assign n2183_o = n2167_o ? n2174_o : n2182_o;
  /* mc8051_tmrctr_rtl.vhd:340:11  */
  assign n2184_o = n2185_o ? n2183_o : s_countl0;
  /* mc8051_tmrctr_rtl.vhd:340:11  */
  assign n2185_o = s_tmr_ctr0_en & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:337:9  */
  assign n2186_o = n2166_o ? reload_i : n2184_o;
  /* mc8051_tmrctr_rtl.vhd:362:17  */
  assign n2188_o = wt_i == 2'b10;
  /* mc8051_tmrctr_rtl.vhd:362:24  */
  assign n2189_o = n2188_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:367:25  */
  assign n2190_o = ~s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:368:29  */
  assign n2192_o = s_count0 == 16'b1111111111111111;
  /* mc8051_tmrctr_rtl.vhd:371:32  */
  assign n2194_o = s_countl0 == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:372:44  */
  assign n2197_o = s_counth0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:371:19  */
  assign n2198_o = n2194_o ? n2197_o : s_counth0;
  /* mc8051_tmrctr_rtl.vhd:368:17  */
  assign n2200_o = n2192_o ? 8'b00000000 : n2198_o;
  /* mc8051_tmrctr_rtl.vhd:377:31  */
  assign n2202_o = s_count0 == 16'b1111111111111111;
  /* mc8051_tmrctr_rtl.vhd:380:34  */
  assign n2204_o = s_countl0 == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:381:46  */
  assign n2207_o = s_counth0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:380:21  */
  assign n2208_o = n2204_o ? n2207_o : s_counth0;
  /* mc8051_tmrctr_rtl.vhd:377:19  */
  assign n2210_o = n2202_o ? 8'b00000000 : n2208_o;
  /* mc8051_tmrctr_rtl.vhd:376:17  */
  assign n2211_o = s_ext_edge0 ? n2210_o : s_counth0;
  /* mc8051_tmrctr_rtl.vhd:367:15  */
  assign n2212_o = n2190_o ? n2200_o : n2211_o;
  /* mc8051_tmrctr_rtl.vhd:365:11  */
  assign n2213_o = n2214_o ? n2212_o : s_counth0;
  /* mc8051_tmrctr_rtl.vhd:365:11  */
  assign n2214_o = s_tmr_ctr0_en & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:362:9  */
  assign n2215_o = n2189_o ? reload_i : n2213_o;
  /* mc8051_tmrctr_rtl.vhd:321:7  */
  assign n2217_o = s_mode0 == 2'b01;
  /* mc8051_tmrctr_rtl.vhd:400:23  */
  assign n2218_o = ~s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:400:51  */
  assign n2219_o = s_ext_edge0 & s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:400:29  */
  assign n2220_o = n2218_o | n2219_o;
  /* mc8051_tmrctr_rtl.vhd:401:26  */
  assign n2221_o = s_count0[7:0];
  /* mc8051_tmrctr_rtl.vhd:401:39  */
  assign n2222_o = {8'b0, n2221_o};  //  uext
  /* mc8051_tmrctr_rtl.vhd:401:39  */
  assign n2224_o = n2222_o == 16'b0000000011111111;
  /* mc8051_tmrctr_rtl.vhd:401:15  */
  assign n2227_o = n2224_o ? 1'b1 : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:400:13  */
  assign n2229_o = n2220_o ? n2227_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:399:11  */
  assign n2231_o = s_count_enable ? n2229_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:398:9  */
  assign n2233_o = s_tmr_ctr0_en ? n2231_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:411:17  */
  assign n2235_o = wt_i == 2'b00;
  /* mc8051_tmrctr_rtl.vhd:411:24  */
  assign n2236_o = n2235_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:416:25  */
  assign n2237_o = ~s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:417:30  */
  assign n2239_o = s_countl0 == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:420:42  */
  assign n2242_o = s_countl0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:417:17  */
  assign n2243_o = n2239_o ? s_counth0 : n2242_o;
  /* mc8051_tmrctr_rtl.vhd:424:32  */
  assign n2245_o = s_countl0 == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:427:44  */
  assign n2248_o = s_countl0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:424:19  */
  assign n2249_o = n2245_o ? s_counth0 : n2248_o;
  /* mc8051_tmrctr_rtl.vhd:423:17  */
  assign n2250_o = s_ext_edge0 ? n2249_o : s_countl0;
  /* mc8051_tmrctr_rtl.vhd:416:15  */
  assign n2251_o = n2237_o ? n2243_o : n2250_o;
  /* mc8051_tmrctr_rtl.vhd:414:11  */
  assign n2252_o = n2253_o ? n2251_o : s_countl0;
  /* mc8051_tmrctr_rtl.vhd:414:11  */
  assign n2253_o = s_tmr_ctr0_en & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:411:9  */
  assign n2254_o = n2236_o ? reload_i : n2252_o;
  /* mc8051_tmrctr_rtl.vhd:436:17  */
  assign n2256_o = wt_i == 2'b10;
  /* mc8051_tmrctr_rtl.vhd:436:24  */
  assign n2257_o = n2256_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:436:9  */
  assign n2258_o = n2257_o ? reload_i : s_counth0;
  /* mc8051_tmrctr_rtl.vhd:395:7  */
  assign n2260_o = s_mode0 == 2'b10;
  /* mc8051_tmrctr_rtl.vhd:449:23  */
  assign n2261_o = ~s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:449:51  */
  assign n2262_o = s_ext_edge0 & s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:449:29  */
  assign n2263_o = n2261_o | n2262_o;
  /* mc8051_tmrctr_rtl.vhd:450:26  */
  assign n2264_o = s_count0[7:0];
  /* mc8051_tmrctr_rtl.vhd:450:39  */
  assign n2265_o = {8'b0, n2264_o};  //  uext
  /* mc8051_tmrctr_rtl.vhd:450:39  */
  assign n2267_o = n2265_o == 16'b0000000011111111;
  /* mc8051_tmrctr_rtl.vhd:450:15  */
  assign n2270_o = n2267_o ? 1'b1 : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:449:13  */
  assign n2272_o = n2263_o ? n2270_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:448:11  */
  assign n2274_o = s_count_enable ? n2272_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:447:9  */
  assign n2276_o = s_tmr_ctr0_en ? n2274_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:460:17  */
  assign n2278_o = wt_i == 2'b00;
  /* mc8051_tmrctr_rtl.vhd:460:24  */
  assign n2279_o = n2278_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:465:25  */
  assign n2280_o = ~s_c_t0;
  /* mc8051_tmrctr_rtl.vhd:466:30  */
  assign n2282_o = s_countl0 == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:469:42  */
  assign n2285_o = s_countl0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:466:17  */
  assign n2287_o = n2282_o ? 8'b00000000 : n2285_o;
  /* mc8051_tmrctr_rtl.vhd:473:32  */
  assign n2289_o = s_countl0 == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:476:44  */
  assign n2292_o = s_countl0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:473:19  */
  assign n2294_o = n2289_o ? 8'b00000000 : n2292_o;
  /* mc8051_tmrctr_rtl.vhd:472:17  */
  assign n2295_o = s_ext_edge0 ? n2294_o : s_countl0;
  /* mc8051_tmrctr_rtl.vhd:465:15  */
  assign n2296_o = n2280_o ? n2287_o : n2295_o;
  /* mc8051_tmrctr_rtl.vhd:463:11  */
  assign n2297_o = n2298_o ? n2296_o : s_countl0;
  /* mc8051_tmrctr_rtl.vhd:463:11  */
  assign n2298_o = s_tmr_ctr0_en & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:460:9  */
  assign n2299_o = n2279_o ? reload_i : n2297_o;
  /* mc8051_tmrctr_rtl.vhd:487:24  */
  assign n2300_o = s_count0[15:8];
  /* mc8051_tmrctr_rtl.vhd:487:38  */
  assign n2302_o = n2300_o == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:487:13  */
  assign n2305_o = n2302_o ? 1'b1 : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:486:11  */
  assign n2307_o = s_count_enable ? n2305_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:485:9  */
  assign n2309_o = tcon_tr1_i ? n2307_o : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:496:17  */
  assign n2311_o = wt_i == 2'b10;
  /* mc8051_tmrctr_rtl.vhd:496:24  */
  assign n2312_o = n2311_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:501:28  */
  assign n2314_o = s_counth0 == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:504:40  */
  assign n2317_o = s_counth0 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:501:15  */
  assign n2319_o = n2314_o ? 8'b00000000 : n2317_o;
  /* mc8051_tmrctr_rtl.vhd:499:11  */
  assign n2320_o = n2321_o ? n2319_o : s_counth0;
  /* mc8051_tmrctr_rtl.vhd:499:11  */
  assign n2321_o = tcon_tr1_i & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:496:9  */
  assign n2322_o = n2312_o ? reload_i : n2320_o;
  /* mc8051_tmrctr_rtl.vhd:444:7  */
  assign n2324_o = s_mode0 == 2'b11;
  assign n2325_o = {n2324_o, n2260_o, n2217_o, n2149_o};
  /* mc8051_tmrctr_rtl.vhd:248:7  */
  always @*
    case (n2325_o)
      4'b1000: n2326_o = n2299_o;
      4'b0100: n2326_o = n2254_o;
      4'b0010: n2326_o = n2186_o;
      4'b0001: n2326_o = n2118_o;
      default: n2326_o = s_countl0;
    endcase
  /* mc8051_tmrctr_rtl.vhd:248:7  */
  always @*
    case (n2325_o)
      4'b1000: n2327_o = n2322_o;
      4'b0100: n2327_o = n2258_o;
      4'b0010: n2327_o = n2215_o;
      4'b0001: n2327_o = n2147_o;
      default: n2327_o = s_counth0;
    endcase
  /* mc8051_tmrctr_rtl.vhd:248:7  */
  always @*
    case (n2325_o)
      4'b1000: n2329_o = n2276_o;
      4'b0100: n2329_o = n2233_o;
      4'b0010: n2329_o = n2163_o;
      4'b0001: n2329_o = n2095_o;
      default: n2329_o = 1'b0;
    endcase
  /* mc8051_tmrctr_rtl.vhd:248:7  */
  always @*
    case (n2325_o)
      4'b1000: n2332_o = n2309_o;
      4'b0100: n2332_o = 1'b0;
      4'b0010: n2332_o = 1'b0;
      4'b0001: n2332_o = 1'b0;
      default: n2332_o = 1'b0;
    endcase
  /* mc8051_tmrctr_rtl.vhd:534:24  */
  assign n2335_o = s_mode0 == 2'b01;
  /* mc8051_tmrctr_rtl.vhd:535:24  */
  assign n2337_o = s_mode0 == 2'b00;
  /* mc8051_tmrctr_rtl.vhd:534:45  */
  assign n2338_o = n2335_o | n2337_o;
  /* mc8051_tmrctr_rtl.vhd:536:24  */
  assign n2340_o = s_mode0 == 2'b10;
  /* mc8051_tmrctr_rtl.vhd:535:45  */
  assign n2341_o = n2338_o | n2340_o;
  /* mc8051_tmrctr_rtl.vhd:537:25  */
  assign n2342_o = ~s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:537:53  */
  assign n2343_o = s_ext_edge1 & s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:537:31  */
  assign n2344_o = n2342_o | n2343_o;
  /* mc8051_tmrctr_rtl.vhd:538:29  */
  assign n2346_o = s_count1 == 16'b1111111100011111;
  /* mc8051_tmrctr_rtl.vhd:538:17  */
  assign n2349_o = n2346_o ? 1'b1 : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:532:9  */
  assign n2350_o = n2353_o ? n2349_o : n2332_o;
  /* mc8051_tmrctr_rtl.vhd:534:13  */
  assign n2351_o = n2341_o & n2344_o;
  /* mc8051_tmrctr_rtl.vhd:533:11  */
  assign n2352_o = s_count_enable & n2351_o;
  /* mc8051_tmrctr_rtl.vhd:532:9  */
  assign n2353_o = s_tmr_ctr1_en & n2352_o;
  /* mc8051_tmrctr_rtl.vhd:551:17  */
  assign n2355_o = wt_i == 2'b01;
  /* mc8051_tmrctr_rtl.vhd:551:24  */
  assign n2356_o = n2355_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:556:25  */
  assign n2357_o = ~s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:557:30  */
  assign n2359_o = s_countl1 == 8'b00011111;
  /* mc8051_tmrctr_rtl.vhd:560:42  */
  assign n2362_o = s_countl1 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:557:17  */
  assign n2364_o = n2359_o ? 8'b00000000 : n2362_o;
  /* mc8051_tmrctr_rtl.vhd:564:32  */
  assign n2366_o = s_countl1 == 8'b00011111;
  /* mc8051_tmrctr_rtl.vhd:567:44  */
  assign n2369_o = s_countl1 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:564:19  */
  assign n2371_o = n2366_o ? 8'b00000000 : n2369_o;
  /* mc8051_tmrctr_rtl.vhd:563:17  */
  assign n2372_o = s_ext_edge1 ? n2371_o : s_countl1;
  /* mc8051_tmrctr_rtl.vhd:556:15  */
  assign n2373_o = n2357_o ? n2364_o : n2372_o;
  /* mc8051_tmrctr_rtl.vhd:554:11  */
  assign n2374_o = n2375_o ? n2373_o : s_countl1;
  /* mc8051_tmrctr_rtl.vhd:554:11  */
  assign n2375_o = s_tmr_ctr1_en & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:551:9  */
  assign n2376_o = n2356_o ? reload_i : n2374_o;
  /* mc8051_tmrctr_rtl.vhd:576:17  */
  assign n2378_o = wt_i == 2'b11;
  /* mc8051_tmrctr_rtl.vhd:576:24  */
  assign n2379_o = n2378_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:581:25  */
  assign n2380_o = ~s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:582:29  */
  assign n2382_o = s_count1 == 16'b1111111100011111;
  /* mc8051_tmrctr_rtl.vhd:585:32  */
  assign n2384_o = s_countl1 == 8'b00011111;
  /* mc8051_tmrctr_rtl.vhd:586:44  */
  assign n2387_o = s_counth1 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:585:19  */
  assign n2388_o = n2384_o ? n2387_o : s_counth1;
  /* mc8051_tmrctr_rtl.vhd:582:17  */
  assign n2390_o = n2382_o ? 8'b00000000 : n2388_o;
  /* mc8051_tmrctr_rtl.vhd:591:31  */
  assign n2392_o = s_count1 == 16'b1111111100011111;
  /* mc8051_tmrctr_rtl.vhd:594:34  */
  assign n2394_o = s_countl1 == 8'b00011111;
  /* mc8051_tmrctr_rtl.vhd:595:46  */
  assign n2397_o = s_counth1 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:594:21  */
  assign n2398_o = n2394_o ? n2397_o : s_counth1;
  /* mc8051_tmrctr_rtl.vhd:591:19  */
  assign n2400_o = n2392_o ? 8'b00000000 : n2398_o;
  /* mc8051_tmrctr_rtl.vhd:590:17  */
  assign n2401_o = s_ext_edge1 ? n2400_o : s_counth1;
  /* mc8051_tmrctr_rtl.vhd:581:15  */
  assign n2402_o = n2380_o ? n2390_o : n2401_o;
  /* mc8051_tmrctr_rtl.vhd:579:11  */
  assign n2403_o = n2404_o ? n2402_o : s_counth1;
  /* mc8051_tmrctr_rtl.vhd:579:11  */
  assign n2404_o = s_tmr_ctr1_en & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:576:9  */
  assign n2405_o = n2379_o ? reload_i : n2403_o;
  /* mc8051_tmrctr_rtl.vhd:529:9  */
  assign n2407_o = s_mode1 == 2'b00;
  /* mc8051_tmrctr_rtl.vhd:612:24  */
  assign n2409_o = s_mode0 == 2'b01;
  /* mc8051_tmrctr_rtl.vhd:613:24  */
  assign n2411_o = s_mode0 == 2'b00;
  /* mc8051_tmrctr_rtl.vhd:612:45  */
  assign n2412_o = n2409_o | n2411_o;
  /* mc8051_tmrctr_rtl.vhd:614:24  */
  assign n2414_o = s_mode0 == 2'b10;
  /* mc8051_tmrctr_rtl.vhd:613:45  */
  assign n2415_o = n2412_o | n2414_o;
  /* mc8051_tmrctr_rtl.vhd:615:25  */
  assign n2416_o = ~s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:615:53  */
  assign n2417_o = s_ext_edge1 & s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:615:31  */
  assign n2418_o = n2416_o | n2417_o;
  /* mc8051_tmrctr_rtl.vhd:616:29  */
  assign n2420_o = s_count1 == 16'b1111111111111111;
  /* mc8051_tmrctr_rtl.vhd:616:17  */
  assign n2423_o = n2420_o ? 1'b1 : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:610:9  */
  assign n2424_o = n2427_o ? n2423_o : n2332_o;
  /* mc8051_tmrctr_rtl.vhd:612:13  */
  assign n2425_o = n2415_o & n2418_o;
  /* mc8051_tmrctr_rtl.vhd:611:11  */
  assign n2426_o = s_count_enable & n2425_o;
  /* mc8051_tmrctr_rtl.vhd:610:9  */
  assign n2427_o = s_tmr_ctr1_en & n2426_o;
  /* mc8051_tmrctr_rtl.vhd:629:17  */
  assign n2429_o = wt_i == 2'b01;
  /* mc8051_tmrctr_rtl.vhd:629:24  */
  assign n2430_o = n2429_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:634:25  */
  assign n2431_o = ~s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:635:29  */
  assign n2433_o = s_count1 == 16'b1111111111111111;
  /* mc8051_tmrctr_rtl.vhd:638:42  */
  assign n2436_o = s_countl1 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:635:17  */
  assign n2438_o = n2433_o ? 8'b00000000 : n2436_o;
  /* mc8051_tmrctr_rtl.vhd:642:31  */
  assign n2440_o = s_count1 == 16'b1111111111111111;
  /* mc8051_tmrctr_rtl.vhd:645:44  */
  assign n2443_o = s_countl1 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:642:19  */
  assign n2445_o = n2440_o ? 8'b00000000 : n2443_o;
  /* mc8051_tmrctr_rtl.vhd:641:17  */
  assign n2446_o = s_ext_edge1 ? n2445_o : s_countl1;
  /* mc8051_tmrctr_rtl.vhd:634:15  */
  assign n2447_o = n2431_o ? n2438_o : n2446_o;
  /* mc8051_tmrctr_rtl.vhd:632:11  */
  assign n2448_o = n2449_o ? n2447_o : s_countl1;
  /* mc8051_tmrctr_rtl.vhd:632:11  */
  assign n2449_o = s_tmr_ctr1_en & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:629:9  */
  assign n2450_o = n2430_o ? reload_i : n2448_o;
  /* mc8051_tmrctr_rtl.vhd:654:17  */
  assign n2452_o = wt_i == 2'b11;
  /* mc8051_tmrctr_rtl.vhd:654:24  */
  assign n2453_o = n2452_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:659:25  */
  assign n2454_o = ~s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:660:29  */
  assign n2456_o = s_count1 == 16'b1111111111111111;
  /* mc8051_tmrctr_rtl.vhd:663:32  */
  assign n2458_o = s_countl1 == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:664:44  */
  assign n2461_o = s_counth1 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:663:19  */
  assign n2462_o = n2458_o ? n2461_o : s_counth1;
  /* mc8051_tmrctr_rtl.vhd:660:17  */
  assign n2464_o = n2456_o ? 8'b00000000 : n2462_o;
  /* mc8051_tmrctr_rtl.vhd:669:31  */
  assign n2466_o = s_count1 == 16'b1111111111111111;
  /* mc8051_tmrctr_rtl.vhd:672:34  */
  assign n2468_o = s_countl1 == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:673:46  */
  assign n2471_o = s_counth1 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:672:21  */
  assign n2472_o = n2468_o ? n2471_o : s_counth1;
  /* mc8051_tmrctr_rtl.vhd:669:19  */
  assign n2474_o = n2466_o ? 8'b00000000 : n2472_o;
  /* mc8051_tmrctr_rtl.vhd:668:17  */
  assign n2475_o = s_ext_edge1 ? n2474_o : s_counth1;
  /* mc8051_tmrctr_rtl.vhd:659:15  */
  assign n2476_o = n2454_o ? n2464_o : n2475_o;
  /* mc8051_tmrctr_rtl.vhd:657:11  */
  assign n2477_o = n2478_o ? n2476_o : s_counth1;
  /* mc8051_tmrctr_rtl.vhd:657:11  */
  assign n2478_o = s_tmr_ctr1_en & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:654:9  */
  assign n2479_o = n2453_o ? reload_i : n2477_o;
  /* mc8051_tmrctr_rtl.vhd:607:9  */
  assign n2481_o = s_mode1 == 2'b01;
  /* mc8051_tmrctr_rtl.vhd:691:24  */
  assign n2483_o = s_mode0 == 2'b01;
  /* mc8051_tmrctr_rtl.vhd:692:24  */
  assign n2485_o = s_mode0 == 2'b00;
  /* mc8051_tmrctr_rtl.vhd:691:45  */
  assign n2486_o = n2483_o | n2485_o;
  /* mc8051_tmrctr_rtl.vhd:693:24  */
  assign n2488_o = s_mode0 == 2'b10;
  /* mc8051_tmrctr_rtl.vhd:692:45  */
  assign n2489_o = n2486_o | n2488_o;
  /* mc8051_tmrctr_rtl.vhd:694:25  */
  assign n2490_o = ~s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:694:53  */
  assign n2491_o = s_ext_edge1 & s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:694:31  */
  assign n2492_o = n2490_o | n2491_o;
  /* mc8051_tmrctr_rtl.vhd:695:28  */
  assign n2493_o = s_count1[7:0];
  /* mc8051_tmrctr_rtl.vhd:695:41  */
  assign n2494_o = {8'b0, n2493_o};  //  uext
  /* mc8051_tmrctr_rtl.vhd:695:41  */
  assign n2496_o = n2494_o == 16'b0000000011111111;
  /* mc8051_tmrctr_rtl.vhd:695:17  */
  assign n2499_o = n2496_o ? 1'b1 : 1'b0;
  /* mc8051_tmrctr_rtl.vhd:689:9  */
  assign n2500_o = n2503_o ? n2499_o : n2332_o;
  /* mc8051_tmrctr_rtl.vhd:691:13  */
  assign n2501_o = n2489_o & n2492_o;
  /* mc8051_tmrctr_rtl.vhd:690:11  */
  assign n2502_o = s_count_enable & n2501_o;
  /* mc8051_tmrctr_rtl.vhd:689:9  */
  assign n2503_o = s_tmr_ctr1_en & n2502_o;
  /* mc8051_tmrctr_rtl.vhd:708:17  */
  assign n2505_o = wt_i == 2'b01;
  /* mc8051_tmrctr_rtl.vhd:708:24  */
  assign n2506_o = n2505_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:713:25  */
  assign n2507_o = ~s_c_t1;
  /* mc8051_tmrctr_rtl.vhd:714:30  */
  assign n2509_o = s_countl1 == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:717:42  */
  assign n2512_o = s_countl1 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:714:17  */
  assign n2513_o = n2509_o ? s_counth1 : n2512_o;
  /* mc8051_tmrctr_rtl.vhd:721:32  */
  assign n2515_o = s_countl1 == 8'b11111111;
  /* mc8051_tmrctr_rtl.vhd:724:44  */
  assign n2518_o = s_countl1 + 8'b00000001;
  /* mc8051_tmrctr_rtl.vhd:721:19  */
  assign n2519_o = n2515_o ? s_counth1 : n2518_o;
  /* mc8051_tmrctr_rtl.vhd:720:17  */
  assign n2520_o = s_ext_edge1 ? n2519_o : s_countl1;
  /* mc8051_tmrctr_rtl.vhd:713:15  */
  assign n2521_o = n2507_o ? n2513_o : n2520_o;
  /* mc8051_tmrctr_rtl.vhd:711:11  */
  assign n2522_o = n2523_o ? n2521_o : s_countl1;
  /* mc8051_tmrctr_rtl.vhd:711:11  */
  assign n2523_o = s_tmr_ctr1_en & s_count_enable;
  /* mc8051_tmrctr_rtl.vhd:708:9  */
  assign n2524_o = n2506_o ? reload_i : n2522_o;
  /* mc8051_tmrctr_rtl.vhd:733:17  */
  assign n2526_o = wt_i == 2'b11;
  /* mc8051_tmrctr_rtl.vhd:733:24  */
  assign n2527_o = n2526_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:733:9  */
  assign n2528_o = n2527_o ? reload_i : s_counth1;
  /* mc8051_tmrctr_rtl.vhd:686:9  */
  assign n2530_o = s_mode1 == 2'b10;
  /* mc8051_tmrctr_rtl.vhd:744:17  */
  assign n2532_o = wt_i == 2'b01;
  /* mc8051_tmrctr_rtl.vhd:744:24  */
  assign n2533_o = n2532_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:744:9  */
  assign n2534_o = n2533_o ? reload_i : s_countl1;
  /* mc8051_tmrctr_rtl.vhd:749:17  */
  assign n2536_o = wt_i == 2'b11;
  /* mc8051_tmrctr_rtl.vhd:749:24  */
  assign n2537_o = n2536_o & wt_en_i;
  /* mc8051_tmrctr_rtl.vhd:749:9  */
  assign n2538_o = n2537_o ? reload_i : s_counth1;
  /* mc8051_tmrctr_rtl.vhd:741:7  */
  assign n2540_o = s_mode1 == 2'b11;
  assign n2541_o = {n2540_o, n2530_o, n2481_o, n2407_o};
  /* mc8051_tmrctr_rtl.vhd:528:7  */
  always @*
    case (n2541_o)
      4'b1000: n2542_o = n2534_o;
      4'b0100: n2542_o = n2524_o;
      4'b0010: n2542_o = n2450_o;
      4'b0001: n2542_o = n2376_o;
      default: n2542_o = s_countl1;
    endcase
  /* mc8051_tmrctr_rtl.vhd:528:7  */
  always @*
    case (n2541_o)
      4'b1000: n2543_o = n2538_o;
      4'b0100: n2543_o = n2528_o;
      4'b0010: n2543_o = n2479_o;
      4'b0001: n2543_o = n2405_o;
      default: n2543_o = s_counth1;
    endcase
  /* mc8051_tmrctr_rtl.vhd:528:7  */
  always @*
    case (n2541_o)
      4'b1000: n2544_o = n2332_o;
      4'b0100: n2544_o = n2500_o;
      4'b0010: n2544_o = n2424_o;
      4'b0001: n2544_o = n2350_o;
      default: n2544_o = n2332_o;
    endcase
  /* mc8051_tmrctr_rtl.vhd:146:9  */
  assign n2564_o = cen ? n2010_o : s_pre_count;
  /* mc8051_tmrctr_rtl.vhd:146:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2565_q <= 4'b0000;
    else
      n2565_q <= n2564_o;
  /* mc8051_tmrctr_rtl.vhd:141:7  */
  assign n2566_o = {s_counth0, s_countl0};
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  assign n2567_o = cen ? n2326_o : s_countl0;
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2568_q <= 8'b00000000;
    else
      n2568_q <= n2567_o;
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  assign n2569_o = cen ? n2327_o : s_counth0;
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2570_q <= 8'b00000000;
    else
      n2570_q <= n2569_o;
  /* mc8051_tmrctr_rtl.vhd:230:5  */
  assign n2571_o = {s_counth1, s_countl1};
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  assign n2572_o = cen ? n2542_o : s_countl1;
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2573_q <= 8'b00000000;
    else
      n2573_q <= n2572_o;
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  assign n2574_o = cen ? n2543_o : s_counth1;
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2575_q <= 8'b00000000;
    else
      n2575_q <= n2574_o;
  /* mc8051_tmrctr_rtl.vhd:230:5  */
  assign n2576_o = {n1972_o, n1973_o};
  assign n2577_o = {n1976_o, n1977_o};
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  assign n2578_o = cen ? n2329_o : s_tf0;
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2579_q <= 1'b0;
    else
      n2579_q <= n2578_o;
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  assign n2580_o = cen ? n2544_o : s_tf1;
  /* mc8051_tmrctr_rtl.vhd:241:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2581_q <= 1'b0;
    else
      n2581_q <= n2580_o;
  /* mc8051_tmrctr_rtl.vhd:178:9  */
  assign n2582_o = cen & n2039_o;
  /* mc8051_tmrctr_rtl.vhd:178:9  */
  assign n2583_o = n2582_o ? t0_i : s_t0ff0;
  /* mc8051_tmrctr_rtl.vhd:178:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2584_q <= 1'b0;
    else
      n2584_q <= n2583_o;
  /* mc8051_tmrctr_rtl.vhd:178:9  */
  assign n2585_o = cen & n2040_o;
  /* mc8051_tmrctr_rtl.vhd:178:9  */
  assign n2586_o = n2585_o ? s_t0ff0 : s_t0ff1;
  /* mc8051_tmrctr_rtl.vhd:178:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2587_q <= 1'b0;
    else
      n2587_q <= n2586_o;
  /* mc8051_tmrctr_rtl.vhd:178:9  */
  assign n2588_o = n2032_o ? s_t0ff1 : s_t0ff2;
  /* mc8051_tmrctr_rtl.vhd:178:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2589_q <= 1'b0;
    else
      n2589_q <= n2588_o;
  /* mc8051_tmrctr_rtl.vhd:202:9  */
  assign n2590_o = cen & n2066_o;
  /* mc8051_tmrctr_rtl.vhd:202:9  */
  assign n2591_o = n2590_o ? t1_i : s_t1ff0;
  /* mc8051_tmrctr_rtl.vhd:202:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2592_q <= 1'b0;
    else
      n2592_q <= n2591_o;
  /* mc8051_tmrctr_rtl.vhd:202:9  */
  assign n2593_o = cen & n2067_o;
  /* mc8051_tmrctr_rtl.vhd:202:9  */
  assign n2594_o = n2593_o ? s_t1ff0 : s_t1ff1;
  /* mc8051_tmrctr_rtl.vhd:202:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2595_q <= 1'b0;
    else
      n2595_q <= n2594_o;
  /* mc8051_tmrctr_rtl.vhd:202:9  */
  assign n2596_o = n2059_o ? s_t1ff1 : s_t1ff2;
  /* mc8051_tmrctr_rtl.vhd:202:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2597_q <= 1'b0;
    else
      n2597_q <= n2596_o;
  /* mc8051_tmrctr_rtl.vhd:146:9  */
  assign n2598_o = cen ? n2014_o : s_int0_sync;
  /* mc8051_tmrctr_rtl.vhd:146:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2599_q <= 2'b00;
    else
      n2599_q <= n2598_o;
  /* mc8051_tmrctr_rtl.vhd:146:9  */
  assign n2600_o = cen ? n2016_o : s_int1_sync;
  /* mc8051_tmrctr_rtl.vhd:146:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n2601_q <= 2'b00;
    else
      n2601_q <= n2600_o;
endmodule

module mc8051_siu
  (input  clk,
   input  cen,
   input  reset,
   input  tf_i,
   input  trans_i,
   input  rxd_i,
   input  [5:0] scon_i,
   input  [7:0] sbuf_i,
   input  smod_i,
   output [7:0] sbuf_o,
   output [2:0] scon_o,
   output rxdwr_o,
   output rxd_o,
   output txd_o);
  wire [5:0] s_rxpre_count;
  wire [5:0] s_txpre_count;
  wire s_m0_shift_en;
  wire s_m2_rxshift_en;
  wire s_m13_rxshift_en;
  wire s_m2_txshift_en;
  wire s_m13_txshift_en;
  wire s_ff0;
  wire s_ff1;
  wire s_tf;
  wire [1:0] s_mode;
  wire s_sm2;
  wire s_detect;
  wire s_ren;
  wire s_rxd_val;
  wire s_txdm0;
  wire s_ri;
  wire s_trans;
  wire s_recv_done;
  wire s_tran_done;
  wire s_rb8;
  wire s_tb8;
  wire [3:0] s_recv_state;
  wire [3:0] s_tran_state;
  wire s_rxd_ff0;
  wire s_rxd_ff1;
  wire s_rxd_ff2;
  wire s_det_ff0;
  wire s_det_ff1;
  wire [10:0] s_tran_sh;
  wire [7:0] s_recv_sh;
  wire [7:0] s_recv_buf;
  wire s_rxm13_ff0;
  wire s_rxm13_ff1;
  wire s_txm13_ff0;
  wire s_txm13_ff1;
  wire n475_o;
  wire n476_o;
  wire n477_o;
  wire n478_o;
  wire n479_o;
  wire n480_o;
  wire n482_o;
  wire n483_o;
  wire n484_o;
  wire n490_o;
  wire n492_o;
  wire n494_o;
  wire n496_o;
  wire n498_o;
  wire n500_o;
  wire n502_o;
  wire [2:0] n503_o;
  reg n504_o;
  wire n506_o;
  wire [3:0] n518_o;
  wire [4:0] n519_o;
  wire n521_o;
  wire n522_o;
  wire [4:0] n525_o;
  wire n527_o;
  wire n528_o;
  wire n530_o;
  wire n531_o;
  wire n532_o;
  wire n533_o;
  wire n534_o;
  wire n537_o;
  wire n538_o;
  wire n539_o;
  wire [4:0] n542_o;
  wire n544_o;
  wire n545_o;
  wire n547_o;
  wire n548_o;
  wire n549_o;
  wire n550_o;
  wire n551_o;
  wire n554_o;
  wire n555_o;
  wire n556_o;
  wire n562_o;
  wire [5:0] n565_o;
  wire n567_o;
  wire [5:0] n569_o;
  wire n571_o;
  wire [5:0] n574_o;
  wire [5:0] n577_o;
  wire [5:0] n578_o;
  wire [5:0] n579_o;
  wire [5:0] n580_o;
  wire [5:0] n582_o;
  wire n584_o;
  wire [5:0] n587_o;
  wire n589_o;
  wire [5:0] n591_o;
  wire n593_o;
  wire [5:0] n596_o;
  wire [5:0] n599_o;
  wire [5:0] n600_o;
  wire [5:0] n601_o;
  wire [5:0] n602_o;
  wire [5:0] n604_o;
  wire [3:0] n605_o;
  wire n607_o;
  wire n610_o;
  wire [4:0] n611_o;
  wire n613_o;
  wire n616_o;
  wire n617_o;
  wire [3:0] n618_o;
  wire n620_o;
  wire n623_o;
  wire [4:0] n624_o;
  wire n626_o;
  wire n629_o;
  wire n630_o;
  wire n651_o;
  wire n652_o;
  wire n653_o;
  wire n656_o;
  wire n657_o;
  wire n658_o;
  wire n659_o;
  wire n660_o;
  wire n661_o;
  wire n667_o;
  wire n668_o;
  wire n669_o;
  wire n670_o;
  wire n671_o;
  wire n672_o;
  wire n673_o;
  wire n674_o;
  wire n676_o;
  wire n678_o;
  wire n679_o;
  wire n680_o;
  wire n681_o;
  wire n682_o;
  wire n683_o;
  wire n684_o;
  wire n685_o;
  wire n686_o;
  wire n687_o;
  wire n689_o;
  wire [1:0] n690_o;
  reg n691_o;
  reg n692_o;
  wire n694_o;
  wire n696_o;
  wire [3:0] n697_o;
  wire n699_o;
  wire [3:0] n700_o;
  wire n702_o;
  wire n703_o;
  wire [3:0] n704_o;
  wire n706_o;
  wire n707_o;
  wire n708_o;
  wire n709_o;
  wire n710_o;
  wire [4:0] n711_o;
  wire n713_o;
  wire [4:0] n714_o;
  wire n716_o;
  wire n717_o;
  wire [4:0] n718_o;
  wire n720_o;
  wire n721_o;
  wire n722_o;
  wire n723_o;
  wire n724_o;
  wire n725_o;
  wire n726_o;
  wire n727_o;
  wire n729_o;
  wire n731_o;
  wire n732_o;
  wire [4:0] n733_o;
  wire n735_o;
  wire [4:0] n736_o;
  wire n738_o;
  wire n739_o;
  wire [4:0] n740_o;
  wire n742_o;
  wire n743_o;
  wire n744_o;
  wire n745_o;
  wire n746_o;
  wire n748_o;
  wire n750_o;
  wire n751_o;
  wire n753_o;
  wire n754_o;
  wire n755_o;
  wire n756_o;
  wire n757_o;
  wire n758_o;
  wire n759_o;
  wire n760_o;
  wire n762_o;
  wire [1:0] n763_o;
  reg n764_o;
  reg n765_o;
  reg n766_o;
  wire n767_o;
  wire n768_o;
  wire n769_o;
  wire n770_o;
  wire n771_o;
  wire n772_o;
  wire n774_o;
  wire n776_o;
  wire n798_o;
  wire n800_o;
  wire n801_o;
  wire n803_o;
  wire n804_o;
  wire n806_o;
  wire n807_o;
  wire n809_o;
  wire n810_o;
  wire n812_o;
  wire n813_o;
  wire n815_o;
  wire n816_o;
  wire n818_o;
  wire n819_o;
  wire n821_o;
  wire n822_o;
  wire n824_o;
  wire n825_o;
  wire n827_o;
  wire n828_o;
  wire n830_o;
  wire n831_o;
  wire n833_o;
  wire n834_o;
  wire n836_o;
  wire n837_o;
  wire n839_o;
  wire n840_o;
  wire n842_o;
  wire n843_o;
  wire [3:0] n844_o;
  wire n846_o;
  wire [3:0] n847_o;
  wire n849_o;
  wire n850_o;
  wire n851_o;
  wire n852_o;
  wire n854_o;
  wire [9:0] n856_o;
  wire n857_o;
  wire n859_o;
  wire [9:0] n861_o;
  wire n862_o;
  wire n864_o;
  wire [9:0] n866_o;
  wire n867_o;
  wire n869_o;
  wire [9:0] n871_o;
  wire n872_o;
  wire n874_o;
  wire [9:0] n876_o;
  wire n877_o;
  wire n879_o;
  wire [9:0] n881_o;
  wire n882_o;
  wire n884_o;
  wire [9:0] n886_o;
  wire n887_o;
  wire n889_o;
  wire [9:0] n891_o;
  wire n892_o;
  wire n894_o;
  wire n896_o;
  wire n899_o;
  wire n901_o;
  wire n903_o;
  wire [10:0] n904_o;
  wire [10:0] n905_o;
  wire [1:0] n908_o;
  wire [7:0] n909_o;
  reg n918_o;
  reg n919_o;
  reg n921_o;
  wire [9:0] n922_o;
  reg [9:0] n923_o;
  wire n924_o;
  reg n925_o;
  reg [1:0] n934_o;
  wire n935_o;
  wire n936_o;
  wire n937_o;
  wire [10:0] n938_o;
  wire [10:0] n939_o;
  wire [1:0] n941_o;
  wire n943_o;
  wire [9:0] n945_o;
  wire n946_o;
  wire n947_o;
  wire [10:0] n948_o;
  wire [10:0] n949_o;
  wire [1:0] n952_o;
  wire n954_o;
  wire [9:0] n956_o;
  wire n957_o;
  wire n958_o;
  wire [10:0] n959_o;
  wire [10:0] n960_o;
  wire [1:0] n963_o;
  wire n965_o;
  wire [9:0] n967_o;
  wire n968_o;
  wire n969_o;
  wire [10:0] n970_o;
  wire [10:0] n971_o;
  wire [1:0] n974_o;
  wire n976_o;
  wire [9:0] n978_o;
  wire n979_o;
  wire n980_o;
  wire [10:0] n981_o;
  wire [10:0] n982_o;
  wire [1:0] n985_o;
  wire n987_o;
  wire [9:0] n989_o;
  wire n990_o;
  wire n991_o;
  wire [10:0] n992_o;
  wire [10:0] n993_o;
  wire [1:0] n996_o;
  wire n998_o;
  wire [9:0] n1000_o;
  wire n1001_o;
  wire n1002_o;
  wire [10:0] n1003_o;
  wire [10:0] n1004_o;
  wire [1:0] n1007_o;
  wire n1009_o;
  wire [9:0] n1011_o;
  wire n1012_o;
  wire n1013_o;
  wire [10:0] n1014_o;
  wire [10:0] n1015_o;
  wire [1:0] n1018_o;
  wire n1020_o;
  wire [9:0] n1022_o;
  wire n1023_o;
  wire n1024_o;
  wire [10:0] n1025_o;
  wire [10:0] n1026_o;
  wire [1:0] n1029_o;
  wire n1031_o;
  wire [9:0] n1033_o;
  wire n1034_o;
  wire n1035_o;
  wire n1037_o;
  wire [10:0] n1038_o;
  wire [10:0] n1039_o;
  wire [1:0] n1042_o;
  wire n1044_o;
  wire n1049_o;
  wire n1051_o;
  wire [10:0] n1052_o;
  wire [10:0] n1053_o;
  wire [1:0] n1056_o;
  wire n1058_o;
  wire n1060_o;
  wire n1061_o;
  wire [1:0] n1063_o;
  wire [8:0] n1064_o;
  reg n1065_o;
  reg n1066_o;
  reg [10:0] n1067_o;
  reg [1:0] n1068_o;
  wire n1070_o;
  wire [9:0] n1072_o;
  wire n1073_o;
  wire n1074_o;
  wire [10:0] n1075_o;
  wire [10:0] n1076_o;
  wire [1:0] n1079_o;
  wire n1081_o;
  wire [9:0] n1083_o;
  wire n1084_o;
  wire n1085_o;
  wire [10:0] n1086_o;
  wire [10:0] n1087_o;
  wire [1:0] n1090_o;
  wire n1092_o;
  wire [9:0] n1094_o;
  wire n1095_o;
  wire n1096_o;
  wire [10:0] n1097_o;
  wire [10:0] n1098_o;
  wire [1:0] n1101_o;
  wire n1103_o;
  wire [9:0] n1105_o;
  wire n1106_o;
  wire n1107_o;
  wire [10:0] n1108_o;
  wire [10:0] n1109_o;
  wire [1:0] n1112_o;
  wire n1114_o;
  wire [9:0] n1116_o;
  wire n1117_o;
  wire n1118_o;
  wire [10:0] n1119_o;
  wire [10:0] n1120_o;
  wire [1:0] n1123_o;
  wire n1125_o;
  wire [9:0] n1127_o;
  wire n1128_o;
  wire n1129_o;
  wire [10:0] n1130_o;
  wire [10:0] n1131_o;
  wire [1:0] n1134_o;
  wire n1136_o;
  wire [9:0] n1138_o;
  wire n1139_o;
  wire n1140_o;
  wire [10:0] n1141_o;
  wire [10:0] n1142_o;
  wire [1:0] n1145_o;
  wire n1147_o;
  wire [9:0] n1149_o;
  wire n1150_o;
  wire n1151_o;
  wire [10:0] n1152_o;
  wire [10:0] n1153_o;
  wire [1:0] n1156_o;
  wire n1158_o;
  wire [9:0] n1160_o;
  wire n1161_o;
  wire n1162_o;
  wire [10:0] n1163_o;
  wire [10:0] n1164_o;
  wire [1:0] n1167_o;
  wire n1169_o;
  wire [9:0] n1171_o;
  wire n1172_o;
  wire n1173_o;
  wire n1175_o;
  wire [10:0] n1176_o;
  wire [10:0] n1177_o;
  wire [1:0] n1180_o;
  wire n1182_o;
  wire n1187_o;
  wire n1189_o;
  wire [10:0] n1190_o;
  wire [10:0] n1191_o;
  wire [1:0] n1194_o;
  wire n1196_o;
  wire n1198_o;
  wire n1199_o;
  wire [1:0] n1201_o;
  wire [9:0] n1202_o;
  reg n1203_o;
  reg n1204_o;
  reg [10:0] n1205_o;
  reg [1:0] n1206_o;
  wire n1208_o;
  wire [9:0] n1210_o;
  wire n1211_o;
  wire n1212_o;
  wire [10:0] n1213_o;
  wire [10:0] n1214_o;
  wire [1:0] n1217_o;
  wire n1219_o;
  wire [9:0] n1221_o;
  wire n1222_o;
  wire n1223_o;
  wire [10:0] n1224_o;
  wire [10:0] n1225_o;
  wire [1:0] n1228_o;
  wire n1230_o;
  wire [9:0] n1232_o;
  wire n1233_o;
  wire n1234_o;
  wire [10:0] n1235_o;
  wire [10:0] n1236_o;
  wire [1:0] n1239_o;
  wire n1241_o;
  wire [9:0] n1243_o;
  wire n1244_o;
  wire n1245_o;
  wire [10:0] n1246_o;
  wire [10:0] n1247_o;
  wire [1:0] n1250_o;
  wire n1252_o;
  wire [9:0] n1254_o;
  wire n1255_o;
  wire n1256_o;
  wire [10:0] n1257_o;
  wire [10:0] n1258_o;
  wire [1:0] n1261_o;
  wire n1263_o;
  wire [9:0] n1265_o;
  wire n1266_o;
  wire n1267_o;
  wire [10:0] n1268_o;
  wire [10:0] n1269_o;
  wire [1:0] n1272_o;
  wire n1274_o;
  wire [9:0] n1276_o;
  wire n1277_o;
  wire n1278_o;
  wire [10:0] n1279_o;
  wire [10:0] n1280_o;
  wire [1:0] n1283_o;
  wire n1285_o;
  wire [9:0] n1287_o;
  wire n1288_o;
  wire n1289_o;
  wire [10:0] n1290_o;
  wire [10:0] n1291_o;
  wire [1:0] n1294_o;
  wire n1296_o;
  wire [9:0] n1298_o;
  wire n1299_o;
  wire n1300_o;
  wire [10:0] n1301_o;
  wire [10:0] n1302_o;
  wire [1:0] n1305_o;
  wire n1307_o;
  wire [9:0] n1309_o;
  wire n1310_o;
  wire n1311_o;
  wire n1313_o;
  wire [10:0] n1314_o;
  wire [10:0] n1315_o;
  wire [1:0] n1318_o;
  wire n1320_o;
  wire n1325_o;
  wire n1327_o;
  wire [10:0] n1328_o;
  wire [10:0] n1329_o;
  wire [1:0] n1332_o;
  wire n1334_o;
  wire n1336_o;
  wire n1337_o;
  wire [1:0] n1339_o;
  wire [9:0] n1340_o;
  reg n1341_o;
  reg n1342_o;
  reg [10:0] n1343_o;
  reg [1:0] n1344_o;
  wire n1346_o;
  wire [3:0] n1347_o;
  reg n1351_o;
  reg n1355_o;
  reg n1356_o;
  reg n1357_o;
  reg [10:0] n1358_o;
  reg [1:0] n1360_o;
  wire [3:0] n1364_o;
  wire n1366_o;
  wire n1368_o;
  wire [1:0] n1369_o;
  reg [3:0] n1371_o;
  wire n1401_o;
  wire n1402_o;
  wire n1404_o;
  wire [1:0] n1407_o;
  wire n1408_o;
  wire [1:0] n1410_o;
  wire n1412_o;
  wire [6:0] n1413_o;
  wire [7:0] n1414_o;
  wire [7:0] n1415_o;
  wire [1:0] n1418_o;
  wire n1420_o;
  wire [6:0] n1421_o;
  wire [7:0] n1422_o;
  wire [7:0] n1423_o;
  wire [1:0] n1426_o;
  wire n1428_o;
  wire [6:0] n1429_o;
  wire [7:0] n1430_o;
  wire [7:0] n1431_o;
  wire [1:0] n1434_o;
  wire n1436_o;
  wire [6:0] n1437_o;
  wire [7:0] n1438_o;
  wire [7:0] n1439_o;
  wire [1:0] n1442_o;
  wire n1444_o;
  wire [6:0] n1445_o;
  wire [7:0] n1446_o;
  wire [7:0] n1447_o;
  wire [1:0] n1450_o;
  wire n1452_o;
  wire [6:0] n1453_o;
  wire [7:0] n1454_o;
  wire [7:0] n1455_o;
  wire [1:0] n1458_o;
  wire n1460_o;
  wire [6:0] n1461_o;
  wire [7:0] n1462_o;
  wire [7:0] n1463_o;
  wire [1:0] n1466_o;
  wire n1468_o;
  wire [6:0] n1469_o;
  wire [6:0] n1470_o;
  wire n1472_o;
  wire [7:0] n1473_o;
  wire [7:0] n1474_o;
  wire [7:0] n1475_o;
  wire [7:0] n1476_o;
  wire [1:0] n1479_o;
  wire n1481_o;
  wire [8:0] n1482_o;
  reg n1483_o;
  reg [7:0] n1484_o;
  reg [7:0] n1485_o;
  reg [1:0] n1487_o;
  wire n1489_o;
  wire n1490_o;
  wire n1492_o;
  wire [7:0] n1494_o;
  wire [1:0] n1497_o;
  wire n1499_o;
  wire n1500_o;
  wire n1501_o;
  wire [6:0] n1502_o;
  wire [7:0] n1503_o;
  wire [7:0] n1504_o;
  wire [1:0] n1507_o;
  wire [1:0] n1510_o;
  wire n1511_o;
  wire [1:0] n1512_o;
  wire n1513_o;
  wire [1:0] n1515_o;
  wire n1517_o;
  wire [6:0] n1518_o;
  wire [7:0] n1519_o;
  wire [7:0] n1520_o;
  wire [1:0] n1523_o;
  wire n1525_o;
  wire [6:0] n1526_o;
  wire [7:0] n1527_o;
  wire [7:0] n1528_o;
  wire [1:0] n1531_o;
  wire n1533_o;
  wire [6:0] n1534_o;
  wire [7:0] n1535_o;
  wire [7:0] n1536_o;
  wire [1:0] n1539_o;
  wire n1541_o;
  wire [6:0] n1542_o;
  wire [7:0] n1543_o;
  wire [7:0] n1544_o;
  wire [1:0] n1547_o;
  wire n1549_o;
  wire [6:0] n1550_o;
  wire [7:0] n1551_o;
  wire [7:0] n1552_o;
  wire [1:0] n1555_o;
  wire n1557_o;
  wire [6:0] n1558_o;
  wire [7:0] n1559_o;
  wire [7:0] n1560_o;
  wire [1:0] n1563_o;
  wire n1565_o;
  wire [6:0] n1566_o;
  wire [7:0] n1567_o;
  wire [7:0] n1568_o;
  wire [1:0] n1571_o;
  wire n1573_o;
  wire [6:0] n1574_o;
  wire [7:0] n1575_o;
  wire [7:0] n1576_o;
  wire [1:0] n1579_o;
  wire n1581_o;
  wire n1582_o;
  wire n1583_o;
  wire n1584_o;
  wire n1585_o;
  wire n1586_o;
  wire n1587_o;
  wire [3:0] n1588_o;
  wire n1590_o;
  wire [6:0] n1591_o;
  wire n1593_o;
  wire n1594_o;
  wire [7:0] n1595_o;
  wire [7:0] n1596_o;
  wire [7:0] n1597_o;
  wire [1:0] n1600_o;
  wire [1:0] n1603_o;
  wire n1604_o;
  wire n1605_o;
  wire n1606_o;
  wire n1607_o;
  wire [1:0] n1608_o;
  wire n1610_o;
  wire [10:0] n1611_o;
  reg n1612_o;
  reg n1613_o;
  reg [7:0] n1614_o;
  reg [7:0] n1615_o;
  reg [1:0] n1617_o;
  wire n1619_o;
  wire n1620_o;
  wire n1622_o;
  wire [7:0] n1624_o;
  wire [1:0] n1627_o;
  wire n1629_o;
  wire n1630_o;
  wire [6:0] n1631_o;
  wire [7:0] n1632_o;
  wire [7:0] n1633_o;
  wire [1:0] n1636_o;
  wire [1:0] n1639_o;
  wire n1640_o;
  wire [1:0] n1641_o;
  wire n1643_o;
  wire [6:0] n1644_o;
  wire [7:0] n1645_o;
  wire [7:0] n1646_o;
  wire [1:0] n1649_o;
  wire n1651_o;
  wire [6:0] n1652_o;
  wire [7:0] n1653_o;
  wire [7:0] n1654_o;
  wire [1:0] n1657_o;
  wire n1659_o;
  wire [6:0] n1660_o;
  wire [7:0] n1661_o;
  wire [7:0] n1662_o;
  wire [1:0] n1665_o;
  wire n1667_o;
  wire [6:0] n1668_o;
  wire [7:0] n1669_o;
  wire [7:0] n1670_o;
  wire [1:0] n1673_o;
  wire n1675_o;
  wire [6:0] n1676_o;
  wire [7:0] n1677_o;
  wire [7:0] n1678_o;
  wire [1:0] n1681_o;
  wire n1683_o;
  wire [6:0] n1684_o;
  wire [7:0] n1685_o;
  wire [7:0] n1686_o;
  wire [1:0] n1689_o;
  wire n1691_o;
  wire [6:0] n1692_o;
  wire [7:0] n1693_o;
  wire [7:0] n1694_o;
  wire [1:0] n1697_o;
  wire n1699_o;
  wire [6:0] n1700_o;
  wire [7:0] n1701_o;
  wire [7:0] n1702_o;
  wire [1:0] n1705_o;
  wire n1707_o;
  wire n1708_o;
  wire n1709_o;
  wire n1710_o;
  wire n1711_o;
  wire n1712_o;
  wire n1713_o;
  wire [6:0] n1714_o;
  wire n1716_o;
  wire n1717_o;
  wire [7:0] n1718_o;
  wire [7:0] n1719_o;
  wire [7:0] n1720_o;
  wire n1721_o;
  wire n1722_o;
  wire n1723_o;
  wire n1724_o;
  wire [1:0] n1727_o;
  wire n1729_o;
  wire [1:0] n1732_o;
  wire n1734_o;
  wire [11:0] n1735_o;
  reg n1736_o;
  reg n1737_o;
  reg [7:0] n1738_o;
  reg [7:0] n1739_o;
  reg [1:0] n1741_o;
  wire n1743_o;
  wire n1744_o;
  wire n1746_o;
  wire [7:0] n1748_o;
  wire [1:0] n1751_o;
  wire n1753_o;
  wire n1754_o;
  wire n1755_o;
  wire [6:0] n1756_o;
  wire [7:0] n1757_o;
  wire [7:0] n1758_o;
  wire [1:0] n1761_o;
  wire [1:0] n1764_o;
  wire n1765_o;
  wire [1:0] n1766_o;
  wire n1767_o;
  wire [1:0] n1769_o;
  wire n1771_o;
  wire [6:0] n1772_o;
  wire [7:0] n1773_o;
  wire [7:0] n1774_o;
  wire [1:0] n1777_o;
  wire n1779_o;
  wire [6:0] n1780_o;
  wire [7:0] n1781_o;
  wire [7:0] n1782_o;
  wire [1:0] n1785_o;
  wire n1787_o;
  wire [6:0] n1788_o;
  wire [7:0] n1789_o;
  wire [7:0] n1790_o;
  wire [1:0] n1793_o;
  wire n1795_o;
  wire [6:0] n1796_o;
  wire [7:0] n1797_o;
  wire [7:0] n1798_o;
  wire [1:0] n1801_o;
  wire n1803_o;
  wire [6:0] n1804_o;
  wire [7:0] n1805_o;
  wire [7:0] n1806_o;
  wire [1:0] n1809_o;
  wire n1811_o;
  wire [6:0] n1812_o;
  wire [7:0] n1813_o;
  wire [7:0] n1814_o;
  wire [1:0] n1817_o;
  wire n1819_o;
  wire [6:0] n1820_o;
  wire [7:0] n1821_o;
  wire [7:0] n1822_o;
  wire [1:0] n1825_o;
  wire n1827_o;
  wire [6:0] n1828_o;
  wire [7:0] n1829_o;
  wire [7:0] n1830_o;
  wire [1:0] n1833_o;
  wire n1835_o;
  wire n1836_o;
  wire n1837_o;
  wire n1838_o;
  wire n1839_o;
  wire n1840_o;
  wire n1841_o;
  wire [6:0] n1842_o;
  wire n1844_o;
  wire n1845_o;
  wire [7:0] n1846_o;
  wire [7:0] n1847_o;
  wire [7:0] n1848_o;
  wire n1849_o;
  wire n1850_o;
  wire n1851_o;
  wire n1852_o;
  wire [1:0] n1855_o;
  wire n1857_o;
  wire [1:0] n1860_o;
  wire n1862_o;
  wire [11:0] n1863_o;
  reg n1864_o;
  reg n1865_o;
  reg [7:0] n1866_o;
  reg [7:0] n1867_o;
  reg [1:0] n1869_o;
  wire n1871_o;
  wire [3:0] n1872_o;
  reg n1873_o;
  reg n1874_o;
  reg [7:0] n1875_o;
  reg [7:0] n1876_o;
  reg [1:0] n1878_o;
  wire [3:0] n1882_o;
  wire n1884_o;
  wire n1886_o;
  wire [1:0] n1887_o;
  reg [3:0] n1889_o;
  wire [5:0] n1912_o;
  reg [5:0] n1913_q;
  wire [5:0] n1914_o;
  reg [5:0] n1915_q;
  wire n1916_o;
  reg n1917_q;
  wire n1918_o;
  reg n1919_q;
  wire [1:0] n1920_o;
  wire n1921_o;
  reg n1922_q;
  wire n1923_o;
  reg n1924_q;
  wire n1925_o;
  reg n1926_q;
  wire n1927_o;
  reg n1928_q;
  wire n1929_o;
  reg n1930_q;
  wire [3:0] n1931_o;
  reg [3:0] n1932_q;
  wire [3:0] n1933_o;
  reg [3:0] n1934_q;
  wire n1935_o;
  reg n1936_q;
  wire n1937_o;
  reg n1938_q;
  wire n1939_o;
  reg n1940_q;
  wire n1941_o;
  reg n1942_q;
  wire n1943_o;
  reg n1944_q;
  wire [10:0] n1945_o;
  reg [10:0] n1946_q;
  wire [7:0] n1947_o;
  reg [7:0] n1948_q;
  wire [7:0] n1949_o;
  reg [7:0] n1950_q;
  wire n1951_o;
  reg n1952_q;
  wire n1953_o;
  reg n1954_q;
  wire n1955_o;
  reg n1956_q;
  wire n1957_o;
  reg n1958_q;
  wire [2:0] n1959_o;
  wire n1960_o;
  reg n1961_q;
  wire n1962_o;
  reg n1963_q;
  assign sbuf_o = s_recv_buf;
  assign scon_o = n1959_o;
  assign rxdwr_o = n1961_q;
  assign rxd_o = n1963_q;
  assign txd_o = s_txdm0;
  /* mc8051_siu_rtl.vhd:375:35  */
  assign s_rxpre_count = n1913_q; // (signal)
  /* mc8051_siu_rtl.vhd:68:10  */
  assign s_txpre_count = n1915_q; // (signal)
  /* mc8051_siu_rtl.vhd:69:10  */
  assign s_m0_shift_en = n522_o; // (signal)
  /* mc8051_siu_rtl.vhd:71:10  */
  assign s_m2_rxshift_en = n534_o; // (signal)
  /* mc8051_siu_rtl.vhd:72:10  */
  assign s_m13_rxshift_en = n539_o; // (signal)
  /* mc8051_siu_rtl.vhd:73:10  */
  assign s_m2_txshift_en = n551_o; // (signal)
  /* mc8051_siu_rtl.vhd:74:10  */
  assign s_m13_txshift_en = n556_o; // (signal)
  /* mc8051_siu_rtl.vhd:75:10  */
  assign s_ff0 = n1917_q; // (signal)
  /* mc8051_siu_rtl.vhd:76:10  */
  assign s_ff1 = n1919_q; // (signal)
  /* mc8051_siu_rtl.vhd:77:10  */
  assign s_tf = n484_o; // (signal)
  /* mc8051_siu_rtl.vhd:78:10  */
  assign s_mode = n1920_o; // (signal)
  /* mc8051_siu_rtl.vhd:79:10  */
  assign s_sm2 = n478_o; // (signal)
  /* mc8051_siu_rtl.vhd:80:10  */
  assign s_detect = n653_o; // (signal)
  /* mc8051_siu_rtl.vhd:81:10  */
  assign s_ren = n477_o; // (signal)
  /* mc8051_siu_rtl.vhd:82:10  */
  assign s_rxd_val = n661_o; // (signal)
  /* mc8051_siu_rtl.vhd:83:10  */
  assign s_txdm0 = n1922_q; // (signal)
  /* mc8051_siu_rtl.vhd:84:10  */
  assign s_ri = n480_o; // (signal)
  /* mc8051_siu_rtl.vhd:85:10  */
  assign s_trans = n1924_q; // (signal)
  /* mc8051_siu_rtl.vhd:86:10  */
  assign s_recv_done = n1926_q; // (signal)
  /* mc8051_siu_rtl.vhd:87:10  */
  assign s_tran_done = n1928_q; // (signal)
  /* mc8051_siu_rtl.vhd:88:10  */
  assign s_rb8 = n1930_q; // (signal)
  /* mc8051_siu_rtl.vhd:89:10  */
  assign s_tb8 = n479_o; // (signal)
  /* mc8051_siu_rtl.vhd:90:10  */
  assign s_recv_state = n1932_q; // (signal)
  /* mc8051_siu_rtl.vhd:91:10  */
  assign s_tran_state = n1934_q; // (signal)
  /* mc8051_siu_rtl.vhd:92:10  */
  assign s_rxd_ff0 = n1936_q; // (signal)
  /* mc8051_siu_rtl.vhd:93:10  */
  assign s_rxd_ff1 = n1938_q; // (signal)
  /* mc8051_siu_rtl.vhd:94:10  */
  assign s_rxd_ff2 = n1940_q; // (signal)
  /* mc8051_siu_rtl.vhd:95:10  */
  assign s_det_ff0 = n1942_q; // (signal)
  /* mc8051_siu_rtl.vhd:96:10  */
  assign s_det_ff1 = n1944_q; // (signal)
  /* mc8051_siu_rtl.vhd:97:10  */
  assign s_tran_sh = n1946_q; // (signal)
  /* mc8051_siu_rtl.vhd:1167:42  */
  assign s_recv_sh = n1948_q; // (signal)
  /* mc8051_siu_rtl.vhd:99:10  */
  assign s_recv_buf = n1950_q; // (signal)
  /* mc8051_siu_rtl.vhd:100:10  */
  assign s_rxm13_ff0 = n1952_q; // (signal)
  /* mc8051_siu_rtl.vhd:101:10  */
  assign s_rxm13_ff1 = n1954_q; // (signal)
  /* mc8051_siu_rtl.vhd:102:10  */
  assign s_txm13_ff0 = n1956_q; // (signal)
  /* mc8051_siu_rtl.vhd:103:10  */
  assign s_txm13_ff1 = n1958_q; // (signal)
  /* mc8051_siu_rtl.vhd:107:22  */
  assign n475_o = scon_i[4];
  /* mc8051_siu_rtl.vhd:108:22  */
  assign n476_o = scon_i[3];
  /* mc8051_siu_rtl.vhd:109:19  */
  assign n477_o = scon_i[1];
  /* mc8051_siu_rtl.vhd:110:19  */
  assign n478_o = scon_i[2];
  /* mc8051_siu_rtl.vhd:111:19  */
  assign n479_o = scon_i[0];
  /* mc8051_siu_rtl.vhd:112:19  */
  assign n480_o = scon_i[5];
  /* mc8051_siu_rtl.vhd:130:43  */
  assign n482_o = ~s_ff1;
  /* mc8051_siu_rtl.vhd:130:33  */
  assign n483_o = s_ff0 & n482_o;
  /* mc8051_siu_rtl.vhd:130:15  */
  assign n484_o = n483_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:150:17  */
  assign n490_o = s_m0_shift_en ? 1'b0 : s_trans;
  /* mc8051_siu_rtl.vhd:149:15  */
  assign n492_o = s_mode == 2'b00;
  /* mc8051_siu_rtl.vhd:154:17  */
  assign n494_o = s_m13_txshift_en ? 1'b0 : s_trans;
  /* mc8051_siu_rtl.vhd:153:15  */
  assign n496_o = s_mode == 2'b01;
  /* mc8051_siu_rtl.vhd:158:17  */
  assign n498_o = s_m2_txshift_en ? 1'b0 : s_trans;
  /* mc8051_siu_rtl.vhd:157:15  */
  assign n500_o = s_mode == 2'b10;
  /* mc8051_siu_rtl.vhd:162:17  */
  assign n502_o = s_m13_txshift_en ? 1'b0 : s_trans;
  /* mc8051_control_struc.vhd:121:3  */
  assign n503_o = {n500_o, n496_o, n492_o};
  /* mc8051_siu_rtl.vhd:148:13  */
  always @*
    case (n503_o)
      3'b100: n504_o = n498_o;
      3'b010: n504_o = n494_o;
      3'b001: n504_o = n490_o;
      default: n504_o = n502_o;
    endcase
  /* mc8051_siu_rtl.vhd:145:11  */
  assign n506_o = trans_i ? 1'b1 : n504_o;
  /* mc8051_siu_rtl.vhd:182:42  */
  assign n518_o = s_txpre_count[3:0];
  /* mc8051_siu_rtl.vhd:182:55  */
  assign n519_o = {1'b0, n518_o};  //  uext
  /* mc8051_siu_rtl.vhd:182:55  */
  assign n521_o = n519_o == 5'b01011;
  /* mc8051_siu_rtl.vhd:182:24  */
  assign n522_o = n521_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:185:45  */
  assign n525_o = s_rxpre_count[4:0];
  /* mc8051_siu_rtl.vhd:185:58  */
  assign n527_o = n525_o == 5'b11111;
  /* mc8051_siu_rtl.vhd:186:32  */
  assign n528_o = n527_o & smod_i;
  /* mc8051_siu_rtl.vhd:187:46  */
  assign n530_o = s_rxpre_count == 6'b111111;
  /* mc8051_siu_rtl.vhd:188:43  */
  assign n531_o = ~smod_i;
  /* mc8051_siu_rtl.vhd:188:32  */
  assign n532_o = n530_o & n531_o;
  /* mc8051_siu_rtl.vhd:186:50  */
  assign n533_o = n528_o | n532_o;
  /* mc8051_siu_rtl.vhd:185:26  */
  assign n534_o = n533_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:190:66  */
  assign n537_o = ~s_rxm13_ff1;
  /* mc8051_siu_rtl.vhd:190:50  */
  assign n538_o = s_rxm13_ff0 & n537_o;
  /* mc8051_siu_rtl.vhd:190:27  */
  assign n539_o = n538_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:193:45  */
  assign n542_o = s_txpre_count[4:0];
  /* mc8051_siu_rtl.vhd:193:58  */
  assign n544_o = n542_o == 5'b11111;
  /* mc8051_siu_rtl.vhd:194:32  */
  assign n545_o = n544_o & smod_i;
  /* mc8051_siu_rtl.vhd:195:46  */
  assign n547_o = s_txpre_count == 6'b111111;
  /* mc8051_siu_rtl.vhd:196:43  */
  assign n548_o = ~smod_i;
  /* mc8051_siu_rtl.vhd:196:32  */
  assign n549_o = n547_o & n548_o;
  /* mc8051_siu_rtl.vhd:194:50  */
  assign n550_o = n545_o | n549_o;
  /* mc8051_siu_rtl.vhd:193:26  */
  assign n551_o = n550_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:198:66  */
  assign n554_o = ~s_txm13_ff1;
  /* mc8051_siu_rtl.vhd:198:50  */
  assign n555_o = s_txm13_ff0 & n554_o;
  /* mc8051_siu_rtl.vhd:198:27  */
  assign n556_o = n555_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:221:22  */
  assign n562_o = s_mode == 2'b00;
  /* mc8051_siu_rtl.vhd:222:46  */
  assign n565_o = s_txpre_count + 6'b000001;
  /* mc8051_siu_rtl.vhd:223:32  */
  assign n567_o = s_txpre_count == 6'b001011;
  /* mc8051_siu_rtl.vhd:223:15  */
  assign n569_o = n567_o ? 6'b000000 : n565_o;
  /* mc8051_siu_rtl.vhd:226:25  */
  assign n571_o = s_mode == 2'b10;
  /* mc8051_siu_rtl.vhd:227:46  */
  assign n574_o = s_txpre_count + 6'b000001;
  /* mc8051_siu_rtl.vhd:230:48  */
  assign n577_o = s_txpre_count + 6'b000001;
  /* mc8051_siu_rtl.vhd:229:15  */
  assign n578_o = s_tf ? n577_o : s_txpre_count;
  /* mc8051_siu_rtl.vhd:226:13  */
  assign n579_o = n571_o ? n574_o : n578_o;
  /* mc8051_siu_rtl.vhd:221:13  */
  assign n580_o = n562_o ? n569_o : n579_o;
  /* mc8051_siu_rtl.vhd:218:11  */
  assign n582_o = trans_i ? 6'b000000 : n580_o;
  /* mc8051_siu_rtl.vhd:238:22  */
  assign n584_o = s_mode == 2'b00;
  /* mc8051_siu_rtl.vhd:239:46  */
  assign n587_o = s_rxpre_count + 6'b000001;
  /* mc8051_siu_rtl.vhd:240:32  */
  assign n589_o = s_rxpre_count == 6'b001011;
  /* mc8051_siu_rtl.vhd:240:15  */
  assign n591_o = n589_o ? 6'b000000 : n587_o;
  /* mc8051_siu_rtl.vhd:243:25  */
  assign n593_o = s_mode == 2'b10;
  /* mc8051_siu_rtl.vhd:244:46  */
  assign n596_o = s_rxpre_count + 6'b000001;
  /* mc8051_siu_rtl.vhd:247:48  */
  assign n599_o = s_rxpre_count + 6'b000001;
  /* mc8051_siu_rtl.vhd:246:15  */
  assign n600_o = s_tf ? n599_o : s_rxpre_count;
  /* mc8051_siu_rtl.vhd:243:13  */
  assign n601_o = n593_o ? n596_o : n600_o;
  /* mc8051_siu_rtl.vhd:238:13  */
  assign n602_o = n584_o ? n591_o : n601_o;
  /* mc8051_siu_rtl.vhd:235:11  */
  assign n604_o = s_detect ? 6'b000000 : n602_o;
  /* mc8051_siu_rtl.vhd:253:29  */
  assign n605_o = s_rxpre_count[3:0];
  /* mc8051_siu_rtl.vhd:253:42  */
  assign n607_o = n605_o == 4'b1111;
  /* mc8051_siu_rtl.vhd:253:13  */
  assign n610_o = n607_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:259:29  */
  assign n611_o = s_rxpre_count[4:0];
  /* mc8051_siu_rtl.vhd:259:42  */
  assign n613_o = n611_o == 5'b11111;
  /* mc8051_siu_rtl.vhd:259:13  */
  assign n616_o = n613_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:252:11  */
  assign n617_o = smod_i ? n610_o : n616_o;
  /* mc8051_siu_rtl.vhd:267:29  */
  assign n618_o = s_txpre_count[3:0];
  /* mc8051_siu_rtl.vhd:267:42  */
  assign n620_o = n618_o == 4'b1111;
  /* mc8051_siu_rtl.vhd:267:13  */
  assign n623_o = n620_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:273:29  */
  assign n624_o = s_txpre_count[4:0];
  /* mc8051_siu_rtl.vhd:273:42  */
  assign n626_o = n624_o == 5'b11111;
  /* mc8051_siu_rtl.vhd:273:13  */
  assign n629_o = n626_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:266:11  */
  assign n630_o = smod_i ? n623_o : n629_o;
  /* mc8051_siu_rtl.vhd:291:34  */
  assign n651_o = ~s_det_ff0;
  /* mc8051_siu_rtl.vhd:291:40  */
  assign n652_o = n651_o & s_det_ff1;
  /* mc8051_siu_rtl.vhd:291:19  */
  assign n653_o = n652_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:292:42  */
  assign n656_o = s_rxd_ff0 & s_rxd_ff1;
  /* mc8051_siu_rtl.vhd:293:42  */
  assign n657_o = s_rxd_ff0 & s_rxd_ff2;
  /* mc8051_siu_rtl.vhd:292:63  */
  assign n658_o = n656_o | n657_o;
  /* mc8051_siu_rtl.vhd:294:42  */
  assign n659_o = s_rxd_ff1 & s_rxd_ff2;
  /* mc8051_siu_rtl.vhd:293:63  */
  assign n660_o = n658_o | n659_o;
  /* mc8051_siu_rtl.vhd:292:20  */
  assign n661_o = n660_o ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:306:25  */
  assign n667_o = s_recv_state == 4'b0000;
  /* mc8051_siu_rtl.vhd:311:19  */
  assign n668_o = s_tf ? rxd_i : s_det_ff0;
  /* mc8051_siu_rtl.vhd:311:19  */
  assign n669_o = s_tf ? s_det_ff0 : s_det_ff1;
  /* mc8051_siu_rtl.vhd:316:35  */
  assign n670_o = s_rxpre_count[0];
  /* mc8051_siu_rtl.vhd:316:19  */
  assign n671_o = n670_o ? rxd_i : s_det_ff0;
  /* mc8051_siu_rtl.vhd:316:19  */
  assign n672_o = n670_o ? s_det_ff0 : s_det_ff1;
  /* mc8051_siu_rtl.vhd:310:17  */
  assign n673_o = smod_i ? n668_o : n671_o;
  /* mc8051_siu_rtl.vhd:310:17  */
  assign n674_o = smod_i ? n669_o : n672_o;
  /* mc8051_siu_rtl.vhd:309:15  */
  assign n676_o = s_mode == 2'b01;
  /* mc8051_siu_rtl.vhd:309:27  */
  assign n678_o = s_mode == 2'b11;
  /* mc8051_siu_rtl.vhd:309:27  */
  assign n679_o = n676_o | n678_o;
  /* mc8051_siu_rtl.vhd:323:35  */
  assign n680_o = s_rxpre_count[0];
  /* mc8051_siu_rtl.vhd:323:19  */
  assign n681_o = n680_o ? rxd_i : s_det_ff0;
  /* mc8051_siu_rtl.vhd:323:19  */
  assign n682_o = n680_o ? s_det_ff0 : s_det_ff1;
  /* mc8051_siu_rtl.vhd:328:35  */
  assign n683_o = s_rxpre_count[1];
  /* mc8051_siu_rtl.vhd:328:19  */
  assign n684_o = n683_o ? rxd_i : s_det_ff0;
  /* mc8051_siu_rtl.vhd:328:19  */
  assign n685_o = n683_o ? s_det_ff0 : s_det_ff1;
  /* mc8051_siu_rtl.vhd:322:17  */
  assign n686_o = smod_i ? n681_o : n684_o;
  /* mc8051_siu_rtl.vhd:322:17  */
  assign n687_o = smod_i ? n682_o : n685_o;
  /* mc8051_siu_rtl.vhd:321:15  */
  assign n689_o = s_mode == 2'b10;
  assign n690_o = {n689_o, n679_o};
  /* mc8051_siu_rtl.vhd:308:13  */
  always @*
    case (n690_o)
      2'b10: n691_o = n686_o;
      2'b01: n691_o = n673_o;
      default: n691_o = s_det_ff0;
    endcase
  /* mc8051_siu_rtl.vhd:308:13  */
  always @*
    case (n690_o)
      2'b10: n692_o = n687_o;
      2'b01: n692_o = n674_o;
      default: n692_o = s_det_ff1;
    endcase
  /* mc8051_siu_rtl.vhd:307:11  */
  assign n694_o = s_ren ? n691_o : 1'b0;
  /* mc8051_siu_rtl.vhd:307:11  */
  assign n696_o = s_ren ? n692_o : 1'b0;
  /* mc8051_siu_rtl.vhd:347:35  */
  assign n697_o = s_rxpre_count[3:0];
  /* mc8051_siu_rtl.vhd:347:48  */
  assign n699_o = n697_o == 4'b0111;
  /* mc8051_siu_rtl.vhd:348:35  */
  assign n700_o = s_rxpre_count[3:0];
  /* mc8051_siu_rtl.vhd:348:48  */
  assign n702_o = n700_o == 4'b1000;
  /* mc8051_siu_rtl.vhd:347:69  */
  assign n703_o = n699_o | n702_o;
  /* mc8051_siu_rtl.vhd:349:35  */
  assign n704_o = s_rxpre_count[3:0];
  /* mc8051_siu_rtl.vhd:349:48  */
  assign n706_o = n704_o == 4'b1001;
  /* mc8051_siu_rtl.vhd:348:69  */
  assign n707_o = n703_o | n706_o;
  /* mc8051_siu_rtl.vhd:347:19  */
  assign n708_o = n707_o ? rxd_i : s_rxd_ff0;
  /* mc8051_siu_rtl.vhd:347:19  */
  assign n709_o = n707_o ? s_rxd_ff0 : s_rxd_ff1;
  /* mc8051_siu_rtl.vhd:347:19  */
  assign n710_o = n707_o ? s_rxd_ff1 : s_rxd_ff2;
  /* mc8051_siu_rtl.vhd:355:35  */
  assign n711_o = s_rxpre_count[4:0];
  /* mc8051_siu_rtl.vhd:355:48  */
  assign n713_o = n711_o == 5'b01110;
  /* mc8051_siu_rtl.vhd:356:35  */
  assign n714_o = s_rxpre_count[4:0];
  /* mc8051_siu_rtl.vhd:356:48  */
  assign n716_o = n714_o == 5'b10000;
  /* mc8051_siu_rtl.vhd:355:70  */
  assign n717_o = n713_o | n716_o;
  /* mc8051_siu_rtl.vhd:357:35  */
  assign n718_o = s_rxpre_count[4:0];
  /* mc8051_siu_rtl.vhd:357:48  */
  assign n720_o = n718_o == 5'b10010;
  /* mc8051_siu_rtl.vhd:356:70  */
  assign n721_o = n717_o | n720_o;
  /* mc8051_siu_rtl.vhd:355:19  */
  assign n722_o = n721_o ? rxd_i : s_rxd_ff0;
  /* mc8051_siu_rtl.vhd:355:19  */
  assign n723_o = n721_o ? s_rxd_ff0 : s_rxd_ff1;
  /* mc8051_siu_rtl.vhd:355:19  */
  assign n724_o = n721_o ? s_rxd_ff1 : s_rxd_ff2;
  /* mc8051_siu_rtl.vhd:346:17  */
  assign n725_o = smod_i ? n708_o : n722_o;
  /* mc8051_siu_rtl.vhd:346:17  */
  assign n726_o = smod_i ? n709_o : n723_o;
  /* mc8051_siu_rtl.vhd:346:17  */
  assign n727_o = smod_i ? n710_o : n724_o;
  /* mc8051_siu_rtl.vhd:345:15  */
  assign n729_o = s_mode == 2'b01;
  /* mc8051_siu_rtl.vhd:345:27  */
  assign n731_o = s_mode == 2'b11;
  /* mc8051_siu_rtl.vhd:345:27  */
  assign n732_o = n729_o | n731_o;
  /* mc8051_siu_rtl.vhd:365:35  */
  assign n733_o = s_rxpre_count[4:0];
  /* mc8051_siu_rtl.vhd:365:48  */
  assign n735_o = n733_o == 5'b01110;
  /* mc8051_siu_rtl.vhd:366:35  */
  assign n736_o = s_rxpre_count[4:0];
  /* mc8051_siu_rtl.vhd:366:48  */
  assign n738_o = n736_o == 5'b10000;
  /* mc8051_siu_rtl.vhd:365:70  */
  assign n739_o = n735_o | n738_o;
  /* mc8051_siu_rtl.vhd:367:35  */
  assign n740_o = s_rxpre_count[4:0];
  /* mc8051_siu_rtl.vhd:367:48  */
  assign n742_o = n740_o == 5'b10010;
  /* mc8051_siu_rtl.vhd:366:70  */
  assign n743_o = n739_o | n742_o;
  /* mc8051_siu_rtl.vhd:365:19  */
  assign n744_o = n743_o ? rxd_i : s_rxd_ff0;
  /* mc8051_siu_rtl.vhd:365:19  */
  assign n745_o = n743_o ? s_rxd_ff0 : s_rxd_ff1;
  /* mc8051_siu_rtl.vhd:365:19  */
  assign n746_o = n743_o ? s_rxd_ff1 : s_rxd_ff2;
  /* mc8051_siu_rtl.vhd:373:48  */
  assign n748_o = s_rxpre_count == 6'b011100;
  /* mc8051_siu_rtl.vhd:374:48  */
  assign n750_o = s_rxpre_count == 6'b100000;
  /* mc8051_siu_rtl.vhd:373:70  */
  assign n751_o = n748_o | n750_o;
  /* mc8051_siu_rtl.vhd:375:48  */
  assign n753_o = s_rxpre_count == 6'b100100;
  /* mc8051_siu_rtl.vhd:374:70  */
  assign n754_o = n751_o | n753_o;
  /* mc8051_siu_rtl.vhd:373:19  */
  assign n755_o = n754_o ? rxd_i : s_rxd_ff0;
  /* mc8051_siu_rtl.vhd:373:19  */
  assign n756_o = n754_o ? s_rxd_ff0 : s_rxd_ff1;
  /* mc8051_siu_rtl.vhd:373:19  */
  assign n757_o = n754_o ? s_rxd_ff1 : s_rxd_ff2;
  /* mc8051_siu_rtl.vhd:364:17  */
  assign n758_o = smod_i ? n744_o : n755_o;
  /* mc8051_siu_rtl.vhd:364:17  */
  assign n759_o = smod_i ? n745_o : n756_o;
  /* mc8051_siu_rtl.vhd:364:17  */
  assign n760_o = smod_i ? n746_o : n757_o;
  /* mc8051_siu_rtl.vhd:363:15  */
  assign n762_o = s_mode == 2'b10;
  assign n763_o = {n762_o, n732_o};
  /* mc8051_siu_rtl.vhd:344:13  */
  always @*
    case (n763_o)
      2'b10: n764_o = n758_o;
      2'b01: n764_o = n725_o;
      default: n764_o = s_rxd_ff0;
    endcase
  /* mc8051_siu_rtl.vhd:344:13  */
  always @*
    case (n763_o)
      2'b10: n765_o = n759_o;
      2'b01: n765_o = n726_o;
      default: n765_o = s_rxd_ff1;
    endcase
  /* mc8051_siu_rtl.vhd:344:13  */
  always @*
    case (n763_o)
      2'b10: n766_o = n760_o;
      2'b01: n766_o = n727_o;
      default: n766_o = s_rxd_ff2;
    endcase
  /* mc8051_siu_rtl.vhd:343:11  */
  assign n767_o = s_ren ? n764_o : s_rxd_ff0;
  /* mc8051_siu_rtl.vhd:343:11  */
  assign n768_o = s_ren ? n765_o : s_rxd_ff1;
  /* mc8051_siu_rtl.vhd:343:11  */
  assign n769_o = s_ren ? n766_o : s_rxd_ff2;
  /* mc8051_siu_rtl.vhd:306:9  */
  assign n770_o = n667_o ? s_rxd_ff0 : n767_o;
  /* mc8051_siu_rtl.vhd:306:9  */
  assign n771_o = n667_o ? s_rxd_ff1 : n768_o;
  /* mc8051_siu_rtl.vhd:306:9  */
  assign n772_o = n667_o ? s_rxd_ff2 : n769_o;
  /* mc8051_siu_rtl.vhd:306:9  */
  assign n774_o = n667_o ? n694_o : 1'b0;
  /* mc8051_siu_rtl.vhd:306:9  */
  assign n776_o = n667_o ? n696_o : 1'b0;
  /* mc8051_siu_rtl.vhd:425:29  */
  assign n798_o = s_tran_state == 4'b0001;
  /* mc8051_siu_rtl.vhd:426:28  */
  assign n800_o = s_tran_state == 4'b0010;
  /* mc8051_siu_rtl.vhd:425:51  */
  assign n801_o = n798_o | n800_o;
  /* mc8051_siu_rtl.vhd:427:28  */
  assign n803_o = s_tran_state == 4'b0011;
  /* mc8051_siu_rtl.vhd:426:50  */
  assign n804_o = n801_o | n803_o;
  /* mc8051_siu_rtl.vhd:428:28  */
  assign n806_o = s_tran_state == 4'b0100;
  /* mc8051_siu_rtl.vhd:427:50  */
  assign n807_o = n804_o | n806_o;
  /* mc8051_siu_rtl.vhd:429:28  */
  assign n809_o = s_tran_state == 4'b0101;
  /* mc8051_siu_rtl.vhd:428:50  */
  assign n810_o = n807_o | n809_o;
  /* mc8051_siu_rtl.vhd:430:28  */
  assign n812_o = s_tran_state == 4'b0110;
  /* mc8051_siu_rtl.vhd:429:50  */
  assign n813_o = n810_o | n812_o;
  /* mc8051_siu_rtl.vhd:431:28  */
  assign n815_o = s_tran_state == 4'b0111;
  /* mc8051_siu_rtl.vhd:430:50  */
  assign n816_o = n813_o | n815_o;
  /* mc8051_siu_rtl.vhd:432:28  */
  assign n818_o = s_tran_state == 4'b1000;
  /* mc8051_siu_rtl.vhd:431:50  */
  assign n819_o = n816_o | n818_o;
  /* mc8051_siu_rtl.vhd:433:28  */
  assign n821_o = s_recv_state == 4'b0001;
  /* mc8051_siu_rtl.vhd:432:50  */
  assign n822_o = n819_o | n821_o;
  /* mc8051_siu_rtl.vhd:434:28  */
  assign n824_o = s_recv_state == 4'b0010;
  /* mc8051_siu_rtl.vhd:433:50  */
  assign n825_o = n822_o | n824_o;
  /* mc8051_siu_rtl.vhd:435:28  */
  assign n827_o = s_recv_state == 4'b0011;
  /* mc8051_siu_rtl.vhd:434:50  */
  assign n828_o = n825_o | n827_o;
  /* mc8051_siu_rtl.vhd:436:28  */
  assign n830_o = s_recv_state == 4'b0100;
  /* mc8051_siu_rtl.vhd:435:50  */
  assign n831_o = n828_o | n830_o;
  /* mc8051_siu_rtl.vhd:437:28  */
  assign n833_o = s_recv_state == 4'b0101;
  /* mc8051_siu_rtl.vhd:436:50  */
  assign n834_o = n831_o | n833_o;
  /* mc8051_siu_rtl.vhd:438:28  */
  assign n836_o = s_recv_state == 4'b0110;
  /* mc8051_siu_rtl.vhd:437:50  */
  assign n837_o = n834_o | n836_o;
  /* mc8051_siu_rtl.vhd:439:28  */
  assign n839_o = s_recv_state == 4'b0111;
  /* mc8051_siu_rtl.vhd:438:50  */
  assign n840_o = n837_o | n839_o;
  /* mc8051_siu_rtl.vhd:440:28  */
  assign n842_o = s_recv_state == 4'b1000;
  /* mc8051_siu_rtl.vhd:439:50  */
  assign n843_o = n840_o | n842_o;
  /* mc8051_siu_rtl.vhd:441:31  */
  assign n844_o = s_txpre_count[3:0];
  /* mc8051_siu_rtl.vhd:441:44  */
  assign n846_o = n844_o == 4'b1110;
  /* mc8051_siu_rtl.vhd:442:30  */
  assign n847_o = s_txpre_count[3:0];
  /* mc8051_siu_rtl.vhd:442:43  */
  assign n849_o = n847_o == 4'b0110;
  /* mc8051_siu_rtl.vhd:441:67  */
  assign n850_o = n846_o | n849_o;
  /* mc8051_siu_rtl.vhd:443:28  */
  assign n851_o = ~s_txdm0;
  /* mc8051_siu_rtl.vhd:441:15  */
  assign n852_o = n850_o ? n851_o : s_txdm0;
  /* mc8051_siu_rtl.vhd:425:13  */
  assign n854_o = n843_o ? n852_o : 1'b1;
  /* mc8051_siu_rtl.vhd:453:53  */
  assign n856_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:455:53  */
  assign n857_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:451:17  */
  assign n859_o = s_tran_state == 4'b0001;
  /* mc8051_siu_rtl.vhd:459:53  */
  assign n861_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:461:53  */
  assign n862_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:457:17  */
  assign n864_o = s_tran_state == 4'b0010;
  /* mc8051_siu_rtl.vhd:465:53  */
  assign n866_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:467:53  */
  assign n867_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:463:17  */
  assign n869_o = s_tran_state == 4'b0011;
  /* mc8051_siu_rtl.vhd:471:53  */
  assign n871_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:473:53  */
  assign n872_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:469:17  */
  assign n874_o = s_tran_state == 4'b0100;
  /* mc8051_siu_rtl.vhd:477:53  */
  assign n876_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:479:53  */
  assign n877_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:475:17  */
  assign n879_o = s_tran_state == 4'b0101;
  /* mc8051_siu_rtl.vhd:483:53  */
  assign n881_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:485:53  */
  assign n882_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:481:17  */
  assign n884_o = s_tran_state == 4'b0110;
  /* mc8051_siu_rtl.vhd:489:53  */
  assign n886_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:491:53  */
  assign n887_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:487:17  */
  assign n889_o = s_tran_state == 4'b0111;
  /* mc8051_siu_rtl.vhd:495:53  */
  assign n891_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:498:53  */
  assign n892_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:493:17  */
  assign n894_o = s_tran_state == 4'b1000;
  /* mc8051_siu_rtl.vhd:508:53  */
  assign n896_o = sbuf_i[0];
  /* mc8051_siu_rtl.vhd:503:19  */
  assign n899_o = s_trans ? 1'b1 : 1'b0;
  /* mc8051_siu_rtl.vhd:503:19  */
  assign n901_o = s_trans ? n896_o : n1963_q;
  /* mc8051_siu_rtl.vhd:503:19  */
  assign n903_o = s_trans ? 1'b0 : s_tran_done;
  assign n904_o = {3'b111, sbuf_i};
  /* mc8051_siu_rtl.vhd:503:19  */
  assign n905_o = s_trans ? n904_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:503:19  */
  assign n908_o = s_trans ? 2'b01 : 2'b00;
  assign n909_o = {n894_o, n889_o, n884_o, n879_o, n874_o, n869_o, n864_o, n859_o};
  /* mc8051_siu_rtl.vhd:450:15  */
  always @*
    case (n909_o)
      8'b10000000: n918_o = 1'b1;
      8'b01000000: n918_o = 1'b1;
      8'b00100000: n918_o = 1'b1;
      8'b00010000: n918_o = 1'b1;
      8'b00001000: n918_o = 1'b1;
      8'b00000100: n918_o = 1'b1;
      8'b00000010: n918_o = 1'b1;
      8'b00000001: n918_o = 1'b1;
      default: n918_o = n899_o;
    endcase
  /* mc8051_siu_rtl.vhd:450:15  */
  always @*
    case (n909_o)
      8'b10000000: n919_o = n892_o;
      8'b01000000: n919_o = n887_o;
      8'b00100000: n919_o = n882_o;
      8'b00010000: n919_o = n877_o;
      8'b00001000: n919_o = n872_o;
      8'b00000100: n919_o = n867_o;
      8'b00000010: n919_o = n862_o;
      8'b00000001: n919_o = n857_o;
      default: n919_o = n901_o;
    endcase
  /* mc8051_siu_rtl.vhd:450:15  */
  always @*
    case (n909_o)
      8'b10000000: n921_o = 1'b1;
      8'b01000000: n921_o = s_tran_done;
      8'b00100000: n921_o = s_tran_done;
      8'b00010000: n921_o = s_tran_done;
      8'b00001000: n921_o = s_tran_done;
      8'b00000100: n921_o = s_tran_done;
      8'b00000010: n921_o = s_tran_done;
      8'b00000001: n921_o = s_tran_done;
      default: n921_o = n903_o;
    endcase
  assign n922_o = n905_o[9:0];
  /* mc8051_siu_rtl.vhd:450:15  */
  always @*
    case (n909_o)
      8'b10000000: n923_o = n891_o;
      8'b01000000: n923_o = n886_o;
      8'b00100000: n923_o = n881_o;
      8'b00010000: n923_o = n876_o;
      8'b00001000: n923_o = n871_o;
      8'b00000100: n923_o = n866_o;
      8'b00000010: n923_o = n861_o;
      8'b00000001: n923_o = n856_o;
      default: n923_o = n922_o;
    endcase
  assign n924_o = n905_o[10];
  /* mc8051_siu_rtl.vhd:450:15  */
  always @*
    case (n909_o)
      8'b10000000: n925_o = 1'b1;
      8'b01000000: n925_o = 1'b1;
      8'b00100000: n925_o = 1'b1;
      8'b00010000: n925_o = 1'b1;
      8'b00001000: n925_o = 1'b1;
      8'b00000100: n925_o = 1'b1;
      8'b00000010: n925_o = 1'b1;
      8'b00000001: n925_o = 1'b1;
      default: n925_o = n924_o;
    endcase
  /* mc8051_siu_rtl.vhd:450:15  */
  always @*
    case (n909_o)
      8'b10000000: n934_o = 2'b10;
      8'b01000000: n934_o = 2'b01;
      8'b00100000: n934_o = 2'b01;
      8'b00010000: n934_o = 2'b01;
      8'b00001000: n934_o = 2'b01;
      8'b00000100: n934_o = 2'b01;
      8'b00000010: n934_o = 2'b01;
      8'b00000001: n934_o = 2'b01;
      default: n934_o = n908_o;
    endcase
  /* mc8051_siu_rtl.vhd:449:13  */
  assign n935_o = s_m0_shift_en ? n918_o : n1961_q;
  /* mc8051_siu_rtl.vhd:449:13  */
  assign n936_o = s_m0_shift_en ? n919_o : n1963_q;
  /* mc8051_siu_rtl.vhd:449:13  */
  assign n937_o = s_m0_shift_en ? n921_o : s_tran_done;
  assign n938_o = {n925_o, n923_o};
  /* mc8051_siu_rtl.vhd:449:13  */
  assign n939_o = s_m0_shift_en ? n938_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:449:13  */
  assign n941_o = s_m0_shift_en ? n934_o : 2'b00;
  /* mc8051_siu_rtl.vhd:423:11  */
  assign n943_o = s_mode == 2'b00;
  /* mc8051_siu_rtl.vhd:523:53  */
  assign n945_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:525:53  */
  assign n946_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:521:17  */
  assign n947_o = s_m13_txshift_en ? n946_o : s_txdm0;
  assign n948_o = {1'b1, n945_o};
  /* mc8051_siu_rtl.vhd:521:17  */
  assign n949_o = s_m13_txshift_en ? n948_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:521:17  */
  assign n952_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:520:15  */
  assign n954_o = s_tran_state == 4'b0001;
  /* mc8051_siu_rtl.vhd:530:53  */
  assign n956_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:532:53  */
  assign n957_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:528:17  */
  assign n958_o = s_m13_txshift_en ? n957_o : s_txdm0;
  assign n959_o = {1'b1, n956_o};
  /* mc8051_siu_rtl.vhd:528:17  */
  assign n960_o = s_m13_txshift_en ? n959_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:528:17  */
  assign n963_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:527:15  */
  assign n965_o = s_tran_state == 4'b0010;
  /* mc8051_siu_rtl.vhd:537:53  */
  assign n967_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:539:53  */
  assign n968_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:535:17  */
  assign n969_o = s_m13_txshift_en ? n968_o : s_txdm0;
  assign n970_o = {1'b1, n967_o};
  /* mc8051_siu_rtl.vhd:535:17  */
  assign n971_o = s_m13_txshift_en ? n970_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:535:17  */
  assign n974_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:534:15  */
  assign n976_o = s_tran_state == 4'b0011;
  /* mc8051_siu_rtl.vhd:544:53  */
  assign n978_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:546:53  */
  assign n979_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:542:17  */
  assign n980_o = s_m13_txshift_en ? n979_o : s_txdm0;
  assign n981_o = {1'b1, n978_o};
  /* mc8051_siu_rtl.vhd:542:17  */
  assign n982_o = s_m13_txshift_en ? n981_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:542:17  */
  assign n985_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:541:15  */
  assign n987_o = s_tran_state == 4'b0100;
  /* mc8051_siu_rtl.vhd:551:53  */
  assign n989_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:553:53  */
  assign n990_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:549:17  */
  assign n991_o = s_m13_txshift_en ? n990_o : s_txdm0;
  assign n992_o = {1'b1, n989_o};
  /* mc8051_siu_rtl.vhd:549:17  */
  assign n993_o = s_m13_txshift_en ? n992_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:549:17  */
  assign n996_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:548:15  */
  assign n998_o = s_tran_state == 4'b0101;
  /* mc8051_siu_rtl.vhd:558:53  */
  assign n1000_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:560:53  */
  assign n1001_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:556:17  */
  assign n1002_o = s_m13_txshift_en ? n1001_o : s_txdm0;
  assign n1003_o = {1'b1, n1000_o};
  /* mc8051_siu_rtl.vhd:556:17  */
  assign n1004_o = s_m13_txshift_en ? n1003_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:556:17  */
  assign n1007_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:555:15  */
  assign n1009_o = s_tran_state == 4'b0110;
  /* mc8051_siu_rtl.vhd:565:53  */
  assign n1011_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:567:53  */
  assign n1012_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:563:17  */
  assign n1013_o = s_m13_txshift_en ? n1012_o : s_txdm0;
  assign n1014_o = {1'b1, n1011_o};
  /* mc8051_siu_rtl.vhd:563:17  */
  assign n1015_o = s_m13_txshift_en ? n1014_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:563:17  */
  assign n1018_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:562:15  */
  assign n1020_o = s_tran_state == 4'b0111;
  /* mc8051_siu_rtl.vhd:572:53  */
  assign n1022_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:574:53  */
  assign n1023_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:570:17  */
  assign n1024_o = s_m13_txshift_en ? n1023_o : s_txdm0;
  assign n1025_o = {1'b1, n1022_o};
  /* mc8051_siu_rtl.vhd:570:17  */
  assign n1026_o = s_m13_txshift_en ? n1025_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:570:17  */
  assign n1029_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:569:15  */
  assign n1031_o = s_tran_state == 4'b1000;
  /* mc8051_siu_rtl.vhd:579:53  */
  assign n1033_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:582:53  */
  assign n1034_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:577:17  */
  assign n1035_o = s_m13_txshift_en ? n1034_o : s_txdm0;
  /* mc8051_siu_rtl.vhd:577:17  */
  assign n1037_o = s_m13_txshift_en ? 1'b1 : s_tran_done;
  assign n1038_o = {1'b1, n1033_o};
  /* mc8051_siu_rtl.vhd:577:17  */
  assign n1039_o = s_m13_txshift_en ? n1038_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:577:17  */
  assign n1042_o = s_m13_txshift_en ? 2'b10 : 2'b00;
  /* mc8051_siu_rtl.vhd:576:15  */
  assign n1044_o = s_tran_state == 4'b1001;
  /* mc8051_siu_rtl.vhd:588:19  */
  assign n1049_o = s_trans ? 1'b0 : 1'b1;
  /* mc8051_siu_rtl.vhd:587:17  */
  assign n1051_o = n1060_o ? 1'b0 : s_tran_done;
  assign n1052_o = {2'b11, sbuf_i, 1'b0};
  /* mc8051_siu_rtl.vhd:587:17  */
  assign n1053_o = n1061_o ? n1052_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:588:19  */
  assign n1056_o = s_trans ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:587:17  */
  assign n1058_o = s_m13_txshift_en ? n1049_o : 1'b1;
  /* mc8051_siu_rtl.vhd:587:17  */
  assign n1060_o = s_m13_txshift_en & s_trans;
  /* mc8051_siu_rtl.vhd:587:17  */
  assign n1061_o = s_m13_txshift_en & s_trans;
  /* mc8051_siu_rtl.vhd:587:17  */
  assign n1063_o = s_m13_txshift_en ? n1056_o : 2'b00;
  assign n1064_o = {n1044_o, n1031_o, n1020_o, n1009_o, n998_o, n987_o, n976_o, n965_o, n954_o};
  /* mc8051_siu_rtl.vhd:519:13  */
  always @*
    case (n1064_o)
      9'b100000000: n1065_o = n1035_o;
      9'b010000000: n1065_o = n1024_o;
      9'b001000000: n1065_o = n1013_o;
      9'b000100000: n1065_o = n1002_o;
      9'b000010000: n1065_o = n991_o;
      9'b000001000: n1065_o = n980_o;
      9'b000000100: n1065_o = n969_o;
      9'b000000010: n1065_o = n958_o;
      9'b000000001: n1065_o = n947_o;
      default: n1065_o = n1058_o;
    endcase
  /* mc8051_siu_rtl.vhd:519:13  */
  always @*
    case (n1064_o)
      9'b100000000: n1066_o = n1037_o;
      9'b010000000: n1066_o = s_tran_done;
      9'b001000000: n1066_o = s_tran_done;
      9'b000100000: n1066_o = s_tran_done;
      9'b000010000: n1066_o = s_tran_done;
      9'b000001000: n1066_o = s_tran_done;
      9'b000000100: n1066_o = s_tran_done;
      9'b000000010: n1066_o = s_tran_done;
      9'b000000001: n1066_o = s_tran_done;
      default: n1066_o = n1051_o;
    endcase
  /* mc8051_siu_rtl.vhd:519:13  */
  always @*
    case (n1064_o)
      9'b100000000: n1067_o = n1039_o;
      9'b010000000: n1067_o = n1026_o;
      9'b001000000: n1067_o = n1015_o;
      9'b000100000: n1067_o = n1004_o;
      9'b000010000: n1067_o = n993_o;
      9'b000001000: n1067_o = n982_o;
      9'b000000100: n1067_o = n971_o;
      9'b000000010: n1067_o = n960_o;
      9'b000000001: n1067_o = n949_o;
      default: n1067_o = n1053_o;
    endcase
  /* mc8051_siu_rtl.vhd:519:13  */
  always @*
    case (n1064_o)
      9'b100000000: n1068_o = n1042_o;
      9'b010000000: n1068_o = n1029_o;
      9'b001000000: n1068_o = n1018_o;
      9'b000100000: n1068_o = n1007_o;
      9'b000010000: n1068_o = n996_o;
      9'b000001000: n1068_o = n985_o;
      9'b000000100: n1068_o = n974_o;
      9'b000000010: n1068_o = n963_o;
      9'b000000001: n1068_o = n952_o;
      default: n1068_o = n1063_o;
    endcase
  /* mc8051_siu_rtl.vhd:516:11  */
  assign n1070_o = s_mode == 2'b01;
  /* mc8051_siu_rtl.vhd:608:53  */
  assign n1072_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:610:53  */
  assign n1073_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:606:17  */
  assign n1074_o = s_m2_txshift_en ? n1073_o : s_txdm0;
  assign n1075_o = {1'b1, n1072_o};
  /* mc8051_siu_rtl.vhd:606:17  */
  assign n1076_o = s_m2_txshift_en ? n1075_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:606:17  */
  assign n1079_o = s_m2_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:605:15  */
  assign n1081_o = s_tran_state == 4'b0001;
  /* mc8051_siu_rtl.vhd:615:53  */
  assign n1083_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:617:53  */
  assign n1084_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:613:17  */
  assign n1085_o = s_m2_txshift_en ? n1084_o : s_txdm0;
  assign n1086_o = {1'b1, n1083_o};
  /* mc8051_siu_rtl.vhd:613:17  */
  assign n1087_o = s_m2_txshift_en ? n1086_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:613:17  */
  assign n1090_o = s_m2_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:612:15  */
  assign n1092_o = s_tran_state == 4'b0010;
  /* mc8051_siu_rtl.vhd:622:53  */
  assign n1094_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:624:53  */
  assign n1095_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:620:17  */
  assign n1096_o = s_m2_txshift_en ? n1095_o : s_txdm0;
  assign n1097_o = {1'b1, n1094_o};
  /* mc8051_siu_rtl.vhd:620:17  */
  assign n1098_o = s_m2_txshift_en ? n1097_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:620:17  */
  assign n1101_o = s_m2_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:619:15  */
  assign n1103_o = s_tran_state == 4'b0011;
  /* mc8051_siu_rtl.vhd:629:53  */
  assign n1105_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:631:53  */
  assign n1106_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:627:17  */
  assign n1107_o = s_m2_txshift_en ? n1106_o : s_txdm0;
  assign n1108_o = {1'b1, n1105_o};
  /* mc8051_siu_rtl.vhd:627:17  */
  assign n1109_o = s_m2_txshift_en ? n1108_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:627:17  */
  assign n1112_o = s_m2_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:626:15  */
  assign n1114_o = s_tran_state == 4'b0100;
  /* mc8051_siu_rtl.vhd:636:53  */
  assign n1116_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:638:53  */
  assign n1117_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:634:17  */
  assign n1118_o = s_m2_txshift_en ? n1117_o : s_txdm0;
  assign n1119_o = {1'b1, n1116_o};
  /* mc8051_siu_rtl.vhd:634:17  */
  assign n1120_o = s_m2_txshift_en ? n1119_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:634:17  */
  assign n1123_o = s_m2_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:633:15  */
  assign n1125_o = s_tran_state == 4'b0101;
  /* mc8051_siu_rtl.vhd:643:53  */
  assign n1127_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:645:53  */
  assign n1128_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:641:17  */
  assign n1129_o = s_m2_txshift_en ? n1128_o : s_txdm0;
  assign n1130_o = {1'b1, n1127_o};
  /* mc8051_siu_rtl.vhd:641:17  */
  assign n1131_o = s_m2_txshift_en ? n1130_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:641:17  */
  assign n1134_o = s_m2_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:640:15  */
  assign n1136_o = s_tran_state == 4'b0110;
  /* mc8051_siu_rtl.vhd:650:53  */
  assign n1138_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:652:53  */
  assign n1139_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:648:17  */
  assign n1140_o = s_m2_txshift_en ? n1139_o : s_txdm0;
  assign n1141_o = {1'b1, n1138_o};
  /* mc8051_siu_rtl.vhd:648:17  */
  assign n1142_o = s_m2_txshift_en ? n1141_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:648:17  */
  assign n1145_o = s_m2_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:647:15  */
  assign n1147_o = s_tran_state == 4'b0111;
  /* mc8051_siu_rtl.vhd:657:53  */
  assign n1149_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:659:53  */
  assign n1150_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:655:17  */
  assign n1151_o = s_m2_txshift_en ? n1150_o : s_txdm0;
  assign n1152_o = {1'b1, n1149_o};
  /* mc8051_siu_rtl.vhd:655:17  */
  assign n1153_o = s_m2_txshift_en ? n1152_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:655:17  */
  assign n1156_o = s_m2_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:654:15  */
  assign n1158_o = s_tran_state == 4'b1000;
  /* mc8051_siu_rtl.vhd:664:53  */
  assign n1160_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:666:53  */
  assign n1161_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:662:17  */
  assign n1162_o = s_m2_txshift_en ? n1161_o : s_txdm0;
  assign n1163_o = {1'b1, n1160_o};
  /* mc8051_siu_rtl.vhd:662:17  */
  assign n1164_o = s_m2_txshift_en ? n1163_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:662:17  */
  assign n1167_o = s_m2_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:661:15  */
  assign n1169_o = s_tran_state == 4'b1001;
  /* mc8051_siu_rtl.vhd:671:53  */
  assign n1171_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:674:53  */
  assign n1172_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:669:17  */
  assign n1173_o = s_m2_txshift_en ? n1172_o : s_txdm0;
  /* mc8051_siu_rtl.vhd:669:17  */
  assign n1175_o = s_m2_txshift_en ? 1'b1 : s_tran_done;
  assign n1176_o = {1'b1, n1171_o};
  /* mc8051_siu_rtl.vhd:669:17  */
  assign n1177_o = s_m2_txshift_en ? n1176_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:669:17  */
  assign n1180_o = s_m2_txshift_en ? 2'b10 : 2'b00;
  /* mc8051_siu_rtl.vhd:668:15  */
  assign n1182_o = s_tran_state == 4'b1010;
  /* mc8051_siu_rtl.vhd:680:19  */
  assign n1187_o = s_trans ? 1'b0 : 1'b1;
  /* mc8051_siu_rtl.vhd:679:17  */
  assign n1189_o = n1198_o ? 1'b0 : s_tran_done;
  assign n1190_o = {1'b1, s_tb8, sbuf_i, 1'b0};
  /* mc8051_siu_rtl.vhd:679:17  */
  assign n1191_o = n1199_o ? n1190_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:680:19  */
  assign n1194_o = s_trans ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:679:17  */
  assign n1196_o = s_m2_txshift_en ? n1187_o : 1'b1;
  /* mc8051_siu_rtl.vhd:679:17  */
  assign n1198_o = s_m2_txshift_en & s_trans;
  /* mc8051_siu_rtl.vhd:679:17  */
  assign n1199_o = s_m2_txshift_en & s_trans;
  /* mc8051_siu_rtl.vhd:679:17  */
  assign n1201_o = s_m2_txshift_en ? n1194_o : 2'b00;
  assign n1202_o = {n1182_o, n1169_o, n1158_o, n1147_o, n1136_o, n1125_o, n1114_o, n1103_o, n1092_o, n1081_o};
  /* mc8051_siu_rtl.vhd:604:13  */
  always @*
    case (n1202_o)
      10'b1000000000: n1203_o = n1173_o;
      10'b0100000000: n1203_o = n1162_o;
      10'b0010000000: n1203_o = n1151_o;
      10'b0001000000: n1203_o = n1140_o;
      10'b0000100000: n1203_o = n1129_o;
      10'b0000010000: n1203_o = n1118_o;
      10'b0000001000: n1203_o = n1107_o;
      10'b0000000100: n1203_o = n1096_o;
      10'b0000000010: n1203_o = n1085_o;
      10'b0000000001: n1203_o = n1074_o;
      default: n1203_o = n1196_o;
    endcase
  /* mc8051_siu_rtl.vhd:604:13  */
  always @*
    case (n1202_o)
      10'b1000000000: n1204_o = n1175_o;
      10'b0100000000: n1204_o = s_tran_done;
      10'b0010000000: n1204_o = s_tran_done;
      10'b0001000000: n1204_o = s_tran_done;
      10'b0000100000: n1204_o = s_tran_done;
      10'b0000010000: n1204_o = s_tran_done;
      10'b0000001000: n1204_o = s_tran_done;
      10'b0000000100: n1204_o = s_tran_done;
      10'b0000000010: n1204_o = s_tran_done;
      10'b0000000001: n1204_o = s_tran_done;
      default: n1204_o = n1189_o;
    endcase
  /* mc8051_siu_rtl.vhd:604:13  */
  always @*
    case (n1202_o)
      10'b1000000000: n1205_o = n1177_o;
      10'b0100000000: n1205_o = n1164_o;
      10'b0010000000: n1205_o = n1153_o;
      10'b0001000000: n1205_o = n1142_o;
      10'b0000100000: n1205_o = n1131_o;
      10'b0000010000: n1205_o = n1120_o;
      10'b0000001000: n1205_o = n1109_o;
      10'b0000000100: n1205_o = n1098_o;
      10'b0000000010: n1205_o = n1087_o;
      10'b0000000001: n1205_o = n1076_o;
      default: n1205_o = n1191_o;
    endcase
  /* mc8051_siu_rtl.vhd:604:13  */
  always @*
    case (n1202_o)
      10'b1000000000: n1206_o = n1180_o;
      10'b0100000000: n1206_o = n1167_o;
      10'b0010000000: n1206_o = n1156_o;
      10'b0001000000: n1206_o = n1145_o;
      10'b0000100000: n1206_o = n1134_o;
      10'b0000010000: n1206_o = n1123_o;
      10'b0000001000: n1206_o = n1112_o;
      10'b0000000100: n1206_o = n1101_o;
      10'b0000000010: n1206_o = n1090_o;
      10'b0000000001: n1206_o = n1079_o;
      default: n1206_o = n1201_o;
    endcase
  /* mc8051_siu_rtl.vhd:601:11  */
  assign n1208_o = s_mode == 2'b10;
  /* mc8051_siu_rtl.vhd:701:53  */
  assign n1210_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:703:53  */
  assign n1211_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:699:17  */
  assign n1212_o = s_m13_txshift_en ? n1211_o : s_txdm0;
  assign n1213_o = {1'b1, n1210_o};
  /* mc8051_siu_rtl.vhd:699:17  */
  assign n1214_o = s_m13_txshift_en ? n1213_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:699:17  */
  assign n1217_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:698:15  */
  assign n1219_o = s_tran_state == 4'b0001;
  /* mc8051_siu_rtl.vhd:708:53  */
  assign n1221_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:710:53  */
  assign n1222_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:706:17  */
  assign n1223_o = s_m13_txshift_en ? n1222_o : s_txdm0;
  assign n1224_o = {1'b1, n1221_o};
  /* mc8051_siu_rtl.vhd:706:17  */
  assign n1225_o = s_m13_txshift_en ? n1224_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:706:17  */
  assign n1228_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:705:15  */
  assign n1230_o = s_tran_state == 4'b0010;
  /* mc8051_siu_rtl.vhd:715:53  */
  assign n1232_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:717:53  */
  assign n1233_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:713:17  */
  assign n1234_o = s_m13_txshift_en ? n1233_o : s_txdm0;
  assign n1235_o = {1'b1, n1232_o};
  /* mc8051_siu_rtl.vhd:713:17  */
  assign n1236_o = s_m13_txshift_en ? n1235_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:713:17  */
  assign n1239_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:712:15  */
  assign n1241_o = s_tran_state == 4'b0011;
  /* mc8051_siu_rtl.vhd:722:53  */
  assign n1243_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:724:53  */
  assign n1244_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:720:17  */
  assign n1245_o = s_m13_txshift_en ? n1244_o : s_txdm0;
  assign n1246_o = {1'b1, n1243_o};
  /* mc8051_siu_rtl.vhd:720:17  */
  assign n1247_o = s_m13_txshift_en ? n1246_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:720:17  */
  assign n1250_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:719:15  */
  assign n1252_o = s_tran_state == 4'b0100;
  /* mc8051_siu_rtl.vhd:729:53  */
  assign n1254_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:731:53  */
  assign n1255_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:727:17  */
  assign n1256_o = s_m13_txshift_en ? n1255_o : s_txdm0;
  assign n1257_o = {1'b1, n1254_o};
  /* mc8051_siu_rtl.vhd:727:17  */
  assign n1258_o = s_m13_txshift_en ? n1257_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:727:17  */
  assign n1261_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:726:15  */
  assign n1263_o = s_tran_state == 4'b0101;
  /* mc8051_siu_rtl.vhd:736:53  */
  assign n1265_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:738:53  */
  assign n1266_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:734:17  */
  assign n1267_o = s_m13_txshift_en ? n1266_o : s_txdm0;
  assign n1268_o = {1'b1, n1265_o};
  /* mc8051_siu_rtl.vhd:734:17  */
  assign n1269_o = s_m13_txshift_en ? n1268_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:734:17  */
  assign n1272_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:733:15  */
  assign n1274_o = s_tran_state == 4'b0110;
  /* mc8051_siu_rtl.vhd:743:53  */
  assign n1276_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:745:53  */
  assign n1277_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:741:17  */
  assign n1278_o = s_m13_txshift_en ? n1277_o : s_txdm0;
  assign n1279_o = {1'b1, n1276_o};
  /* mc8051_siu_rtl.vhd:741:17  */
  assign n1280_o = s_m13_txshift_en ? n1279_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:741:17  */
  assign n1283_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:740:15  */
  assign n1285_o = s_tran_state == 4'b0111;
  /* mc8051_siu_rtl.vhd:750:53  */
  assign n1287_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:752:53  */
  assign n1288_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:748:17  */
  assign n1289_o = s_m13_txshift_en ? n1288_o : s_txdm0;
  assign n1290_o = {1'b1, n1287_o};
  /* mc8051_siu_rtl.vhd:748:17  */
  assign n1291_o = s_m13_txshift_en ? n1290_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:748:17  */
  assign n1294_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:747:15  */
  assign n1296_o = s_tran_state == 4'b1000;
  /* mc8051_siu_rtl.vhd:757:53  */
  assign n1298_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:759:53  */
  assign n1299_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:755:17  */
  assign n1300_o = s_m13_txshift_en ? n1299_o : s_txdm0;
  assign n1301_o = {1'b1, n1298_o};
  /* mc8051_siu_rtl.vhd:755:17  */
  assign n1302_o = s_m13_txshift_en ? n1301_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:755:17  */
  assign n1305_o = s_m13_txshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:754:15  */
  assign n1307_o = s_tran_state == 4'b1001;
  /* mc8051_siu_rtl.vhd:764:53  */
  assign n1309_o = s_tran_sh[10:1];
  /* mc8051_siu_rtl.vhd:767:53  */
  assign n1310_o = s_tran_sh[1];
  /* mc8051_siu_rtl.vhd:762:17  */
  assign n1311_o = s_m13_txshift_en ? n1310_o : s_txdm0;
  /* mc8051_siu_rtl.vhd:762:17  */
  assign n1313_o = s_m13_txshift_en ? 1'b1 : s_tran_done;
  assign n1314_o = {1'b1, n1309_o};
  /* mc8051_siu_rtl.vhd:762:17  */
  assign n1315_o = s_m13_txshift_en ? n1314_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:762:17  */
  assign n1318_o = s_m13_txshift_en ? 2'b10 : 2'b00;
  /* mc8051_siu_rtl.vhd:761:15  */
  assign n1320_o = s_tran_state == 4'b1010;
  /* mc8051_siu_rtl.vhd:773:19  */
  assign n1325_o = s_trans ? 1'b0 : 1'b1;
  /* mc8051_siu_rtl.vhd:772:17  */
  assign n1327_o = n1336_o ? 1'b0 : s_tran_done;
  assign n1328_o = {1'b1, s_tb8, sbuf_i, 1'b0};
  /* mc8051_siu_rtl.vhd:772:17  */
  assign n1329_o = n1337_o ? n1328_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:773:19  */
  assign n1332_o = s_trans ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:772:17  */
  assign n1334_o = s_m13_txshift_en ? n1325_o : 1'b1;
  /* mc8051_siu_rtl.vhd:772:17  */
  assign n1336_o = s_m13_txshift_en & s_trans;
  /* mc8051_siu_rtl.vhd:772:17  */
  assign n1337_o = s_m13_txshift_en & s_trans;
  /* mc8051_siu_rtl.vhd:772:17  */
  assign n1339_o = s_m13_txshift_en ? n1332_o : 2'b00;
  assign n1340_o = {n1320_o, n1307_o, n1296_o, n1285_o, n1274_o, n1263_o, n1252_o, n1241_o, n1230_o, n1219_o};
  /* mc8051_siu_rtl.vhd:697:13  */
  always @*
    case (n1340_o)
      10'b1000000000: n1341_o = n1311_o;
      10'b0100000000: n1341_o = n1300_o;
      10'b0010000000: n1341_o = n1289_o;
      10'b0001000000: n1341_o = n1278_o;
      10'b0000100000: n1341_o = n1267_o;
      10'b0000010000: n1341_o = n1256_o;
      10'b0000001000: n1341_o = n1245_o;
      10'b0000000100: n1341_o = n1234_o;
      10'b0000000010: n1341_o = n1223_o;
      10'b0000000001: n1341_o = n1212_o;
      default: n1341_o = n1334_o;
    endcase
  /* mc8051_siu_rtl.vhd:697:13  */
  always @*
    case (n1340_o)
      10'b1000000000: n1342_o = n1313_o;
      10'b0100000000: n1342_o = s_tran_done;
      10'b0010000000: n1342_o = s_tran_done;
      10'b0001000000: n1342_o = s_tran_done;
      10'b0000100000: n1342_o = s_tran_done;
      10'b0000010000: n1342_o = s_tran_done;
      10'b0000001000: n1342_o = s_tran_done;
      10'b0000000100: n1342_o = s_tran_done;
      10'b0000000010: n1342_o = s_tran_done;
      10'b0000000001: n1342_o = s_tran_done;
      default: n1342_o = n1327_o;
    endcase
  /* mc8051_siu_rtl.vhd:697:13  */
  always @*
    case (n1340_o)
      10'b1000000000: n1343_o = n1315_o;
      10'b0100000000: n1343_o = n1302_o;
      10'b0010000000: n1343_o = n1291_o;
      10'b0001000000: n1343_o = n1280_o;
      10'b0000100000: n1343_o = n1269_o;
      10'b0000010000: n1343_o = n1258_o;
      10'b0000001000: n1343_o = n1247_o;
      10'b0000000100: n1343_o = n1236_o;
      10'b0000000010: n1343_o = n1225_o;
      10'b0000000001: n1343_o = n1214_o;
      default: n1343_o = n1329_o;
    endcase
  /* mc8051_siu_rtl.vhd:697:13  */
  always @*
    case (n1340_o)
      10'b1000000000: n1344_o = n1318_o;
      10'b0100000000: n1344_o = n1305_o;
      10'b0010000000: n1344_o = n1294_o;
      10'b0001000000: n1344_o = n1283_o;
      10'b0000100000: n1344_o = n1272_o;
      10'b0000010000: n1344_o = n1261_o;
      10'b0000001000: n1344_o = n1250_o;
      10'b0000000100: n1344_o = n1239_o;
      10'b0000000010: n1344_o = n1228_o;
      10'b0000000001: n1344_o = n1217_o;
      default: n1344_o = n1339_o;
    endcase
  /* mc8051_siu_rtl.vhd:694:11  */
  assign n1346_o = s_mode == 2'b11;
  assign n1347_o = {n1346_o, n1208_o, n1070_o, n943_o};
  /* mc8051_siu_rtl.vhd:419:9  */
  always @*
    case (n1347_o)
      4'b1000: n1351_o = 1'b0;
      4'b0100: n1351_o = 1'b0;
      4'b0010: n1351_o = 1'b0;
      4'b0001: n1351_o = n935_o;
      default: n1351_o = n1961_q;
    endcase
  /* mc8051_siu_rtl.vhd:419:9  */
  always @*
    case (n1347_o)
      4'b1000: n1355_o = 1'b0;
      4'b0100: n1355_o = 1'b0;
      4'b0010: n1355_o = 1'b0;
      4'b0001: n1355_o = n936_o;
      default: n1355_o = n1963_q;
    endcase
  /* mc8051_siu_rtl.vhd:419:9  */
  always @*
    case (n1347_o)
      4'b1000: n1356_o = n1341_o;
      4'b0100: n1356_o = n1203_o;
      4'b0010: n1356_o = n1065_o;
      4'b0001: n1356_o = n854_o;
      default: n1356_o = s_txdm0;
    endcase
  /* mc8051_siu_rtl.vhd:419:9  */
  always @*
    case (n1347_o)
      4'b1000: n1357_o = n1342_o;
      4'b0100: n1357_o = n1204_o;
      4'b0010: n1357_o = n1066_o;
      4'b0001: n1357_o = n937_o;
      default: n1357_o = s_tran_done;
    endcase
  /* mc8051_siu_rtl.vhd:419:9  */
  always @*
    case (n1347_o)
      4'b1000: n1358_o = n1343_o;
      4'b0100: n1358_o = n1205_o;
      4'b0010: n1358_o = n1067_o;
      4'b0001: n1358_o = n939_o;
      default: n1358_o = s_tran_sh;
    endcase
  /* mc8051_siu_rtl.vhd:419:9  */
  always @*
    case (n1347_o)
      4'b1000: n1360_o = n1344_o;
      4'b0100: n1360_o = n1206_o;
      4'b0010: n1360_o = n1068_o;
      4'b0001: n1360_o = n941_o;
      default: n1360_o = 2'b00;
    endcase
  /* mc8051_siu_rtl.vhd:791:42  */
  assign n1364_o = s_tran_state + 4'b0001;
  /* mc8051_siu_rtl.vhd:790:11  */
  assign n1366_o = n1360_o == 2'b01;
  /* mc8051_siu_rtl.vhd:792:11  */
  assign n1368_o = n1360_o == 2'b10;
  assign n1369_o = {n1368_o, n1366_o};
  /* mc8051_siu_rtl.vhd:789:9  */
  always @*
    case (n1369_o)
      2'b10: n1371_o = 4'b0000;
      2'b01: n1371_o = n1364_o;
      default: n1371_o = s_tran_state;
    endcase
  /* mc8051_siu_rtl.vhd:830:39  */
  assign n1401_o = ~s_ri;
  /* mc8051_siu_rtl.vhd:830:30  */
  assign n1402_o = s_ren & n1401_o;
  /* mc8051_siu_rtl.vhd:830:15  */
  assign n1404_o = n1408_o ? 1'b0 : s_recv_done;
  /* mc8051_siu_rtl.vhd:831:17  */
  assign n1407_o = s_m0_shift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:830:15  */
  assign n1408_o = n1402_o & s_m0_shift_en;
  /* mc8051_siu_rtl.vhd:830:15  */
  assign n1410_o = n1402_o ? n1407_o : 2'b00;
  /* mc8051_siu_rtl.vhd:828:13  */
  assign n1412_o = s_recv_state == 4'b0000;
  /* mc8051_siu_rtl.vhd:839:51  */
  assign n1413_o = s_recv_sh[7:1];
  assign n1414_o = {rxd_i, n1413_o};
  /* mc8051_siu_rtl.vhd:837:15  */
  assign n1415_o = s_m0_shift_en ? n1414_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:837:15  */
  assign n1418_o = s_m0_shift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:836:13  */
  assign n1420_o = s_recv_state == 4'b0001;
  /* mc8051_siu_rtl.vhd:845:51  */
  assign n1421_o = s_recv_sh[7:1];
  assign n1422_o = {rxd_i, n1421_o};
  /* mc8051_siu_rtl.vhd:843:15  */
  assign n1423_o = s_m0_shift_en ? n1422_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:843:15  */
  assign n1426_o = s_m0_shift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:842:13  */
  assign n1428_o = s_recv_state == 4'b0010;
  /* mc8051_siu_rtl.vhd:851:51  */
  assign n1429_o = s_recv_sh[7:1];
  assign n1430_o = {rxd_i, n1429_o};
  /* mc8051_siu_rtl.vhd:849:15  */
  assign n1431_o = s_m0_shift_en ? n1430_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:849:15  */
  assign n1434_o = s_m0_shift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:848:13  */
  assign n1436_o = s_recv_state == 4'b0011;
  /* mc8051_siu_rtl.vhd:857:51  */
  assign n1437_o = s_recv_sh[7:1];
  assign n1438_o = {rxd_i, n1437_o};
  /* mc8051_siu_rtl.vhd:855:15  */
  assign n1439_o = s_m0_shift_en ? n1438_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:855:15  */
  assign n1442_o = s_m0_shift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:854:13  */
  assign n1444_o = s_recv_state == 4'b0100;
  /* mc8051_siu_rtl.vhd:863:51  */
  assign n1445_o = s_recv_sh[7:1];
  assign n1446_o = {rxd_i, n1445_o};
  /* mc8051_siu_rtl.vhd:861:15  */
  assign n1447_o = s_m0_shift_en ? n1446_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:861:15  */
  assign n1450_o = s_m0_shift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:860:13  */
  assign n1452_o = s_recv_state == 4'b0101;
  /* mc8051_siu_rtl.vhd:869:51  */
  assign n1453_o = s_recv_sh[7:1];
  assign n1454_o = {rxd_i, n1453_o};
  /* mc8051_siu_rtl.vhd:867:15  */
  assign n1455_o = s_m0_shift_en ? n1454_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:867:15  */
  assign n1458_o = s_m0_shift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:866:13  */
  assign n1460_o = s_recv_state == 4'b0110;
  /* mc8051_siu_rtl.vhd:875:51  */
  assign n1461_o = s_recv_sh[7:1];
  assign n1462_o = {rxd_i, n1461_o};
  /* mc8051_siu_rtl.vhd:873:15  */
  assign n1463_o = s_m0_shift_en ? n1462_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:873:15  */
  assign n1466_o = s_m0_shift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:872:13  */
  assign n1468_o = s_recv_state == 4'b0111;
  /* mc8051_siu_rtl.vhd:881:51  */
  assign n1469_o = s_recv_sh[7:1];
  /* mc8051_siu_rtl.vhd:884:52  */
  assign n1470_o = s_recv_sh[7:1];
  /* mc8051_siu_rtl.vhd:879:15  */
  assign n1472_o = s_m0_shift_en ? 1'b1 : s_recv_done;
  assign n1473_o = {rxd_i, n1469_o};
  /* mc8051_siu_rtl.vhd:879:15  */
  assign n1474_o = s_m0_shift_en ? n1473_o : s_recv_sh;
  assign n1475_o = {rxd_i, n1470_o};
  /* mc8051_siu_rtl.vhd:879:15  */
  assign n1476_o = s_m0_shift_en ? n1475_o : s_recv_buf;
  /* mc8051_siu_rtl.vhd:879:15  */
  assign n1479_o = s_m0_shift_en ? 2'b10 : 2'b00;
  /* mc8051_siu_rtl.vhd:878:13  */
  assign n1481_o = s_recv_state == 4'b1000;
  assign n1482_o = {n1481_o, n1468_o, n1460_o, n1452_o, n1444_o, n1436_o, n1428_o, n1420_o, n1412_o};
  /* mc8051_siu_rtl.vhd:827:13  */
  always @*
    case (n1482_o)
      9'b100000000: n1483_o = n1472_o;
      9'b010000000: n1483_o = s_recv_done;
      9'b001000000: n1483_o = s_recv_done;
      9'b000100000: n1483_o = s_recv_done;
      9'b000010000: n1483_o = s_recv_done;
      9'b000001000: n1483_o = s_recv_done;
      9'b000000100: n1483_o = s_recv_done;
      9'b000000010: n1483_o = s_recv_done;
      9'b000000001: n1483_o = n1404_o;
      default: n1483_o = s_recv_done;
    endcase
  /* mc8051_siu_rtl.vhd:827:13  */
  always @*
    case (n1482_o)
      9'b100000000: n1484_o = n1474_o;
      9'b010000000: n1484_o = n1463_o;
      9'b001000000: n1484_o = n1455_o;
      9'b000100000: n1484_o = n1447_o;
      9'b000010000: n1484_o = n1439_o;
      9'b000001000: n1484_o = n1431_o;
      9'b000000100: n1484_o = n1423_o;
      9'b000000010: n1484_o = n1415_o;
      9'b000000001: n1484_o = s_recv_sh;
      default: n1484_o = s_recv_sh;
    endcase
  /* mc8051_siu_rtl.vhd:827:13  */
  always @*
    case (n1482_o)
      9'b100000000: n1485_o = n1476_o;
      9'b010000000: n1485_o = s_recv_buf;
      9'b001000000: n1485_o = s_recv_buf;
      9'b000100000: n1485_o = s_recv_buf;
      9'b000010000: n1485_o = s_recv_buf;
      9'b000001000: n1485_o = s_recv_buf;
      9'b000000100: n1485_o = s_recv_buf;
      9'b000000010: n1485_o = s_recv_buf;
      9'b000000001: n1485_o = s_recv_buf;
      default: n1485_o = s_recv_buf;
    endcase
  /* mc8051_siu_rtl.vhd:827:13  */
  always @*
    case (n1482_o)
      9'b100000000: n1487_o = n1479_o;
      9'b010000000: n1487_o = n1466_o;
      9'b001000000: n1487_o = n1458_o;
      9'b000100000: n1487_o = n1450_o;
      9'b000010000: n1487_o = n1442_o;
      9'b000001000: n1487_o = n1434_o;
      9'b000000100: n1487_o = n1426_o;
      9'b000000010: n1487_o = n1418_o;
      9'b000000001: n1487_o = n1410_o;
      default: n1487_o = 2'b10;
    endcase
  /* mc8051_siu_rtl.vhd:826:11  */
  assign n1489_o = s_mode == 2'b00;
  /* mc8051_siu_rtl.vhd:897:30  */
  assign n1490_o = s_ren & s_detect;
  /* mc8051_siu_rtl.vhd:897:15  */
  assign n1492_o = n1490_o ? 1'b0 : s_recv_done;
  /* mc8051_siu_rtl.vhd:897:15  */
  assign n1494_o = n1490_o ? 8'b00000000 : s_recv_sh;
  /* mc8051_siu_rtl.vhd:897:15  */
  assign n1497_o = n1490_o ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:896:13  */
  assign n1499_o = s_recv_state == 4'b0000;
  /* mc8051_siu_rtl.vhd:903:27  */
  assign n1500_o = ~s_detect;
  /* mc8051_siu_rtl.vhd:904:30  */
  assign n1501_o = ~s_rxd_val;
  /* mc8051_siu_rtl.vhd:907:55  */
  assign n1502_o = s_recv_sh[7:1];
  assign n1503_o = {s_rxd_val, n1502_o};
  /* mc8051_siu_rtl.vhd:903:15  */
  assign n1504_o = n1513_o ? n1503_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:905:19  */
  assign n1507_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:911:19  */
  assign n1510_o = s_m13_rxshift_en ? 2'b10 : 2'b00;
  /* mc8051_siu_rtl.vhd:904:17  */
  assign n1511_o = n1501_o & s_m13_rxshift_en;
  /* mc8051_siu_rtl.vhd:904:17  */
  assign n1512_o = n1501_o ? n1507_o : n1510_o;
  /* mc8051_siu_rtl.vhd:903:15  */
  assign n1513_o = n1500_o & n1511_o;
  /* mc8051_siu_rtl.vhd:903:15  */
  assign n1515_o = n1500_o ? n1512_o : 2'b00;
  /* mc8051_siu_rtl.vhd:902:13  */
  assign n1517_o = s_recv_state == 4'b0001;
  /* mc8051_siu_rtl.vhd:919:51  */
  assign n1518_o = s_recv_sh[7:1];
  assign n1519_o = {s_rxd_val, n1518_o};
  /* mc8051_siu_rtl.vhd:917:15  */
  assign n1520_o = s_m13_rxshift_en ? n1519_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:917:15  */
  assign n1523_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:916:13  */
  assign n1525_o = s_recv_state == 4'b0010;
  /* mc8051_siu_rtl.vhd:925:51  */
  assign n1526_o = s_recv_sh[7:1];
  assign n1527_o = {s_rxd_val, n1526_o};
  /* mc8051_siu_rtl.vhd:923:15  */
  assign n1528_o = s_m13_rxshift_en ? n1527_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:923:15  */
  assign n1531_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:922:13  */
  assign n1533_o = s_recv_state == 4'b0011;
  /* mc8051_siu_rtl.vhd:931:51  */
  assign n1534_o = s_recv_sh[7:1];
  assign n1535_o = {s_rxd_val, n1534_o};
  /* mc8051_siu_rtl.vhd:929:15  */
  assign n1536_o = s_m13_rxshift_en ? n1535_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:929:15  */
  assign n1539_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:928:13  */
  assign n1541_o = s_recv_state == 4'b0100;
  /* mc8051_siu_rtl.vhd:937:51  */
  assign n1542_o = s_recv_sh[7:1];
  assign n1543_o = {s_rxd_val, n1542_o};
  /* mc8051_siu_rtl.vhd:935:15  */
  assign n1544_o = s_m13_rxshift_en ? n1543_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:935:15  */
  assign n1547_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:934:13  */
  assign n1549_o = s_recv_state == 4'b0101;
  /* mc8051_siu_rtl.vhd:943:51  */
  assign n1550_o = s_recv_sh[7:1];
  assign n1551_o = {s_rxd_val, n1550_o};
  /* mc8051_siu_rtl.vhd:941:15  */
  assign n1552_o = s_m13_rxshift_en ? n1551_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:941:15  */
  assign n1555_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:940:13  */
  assign n1557_o = s_recv_state == 4'b0110;
  /* mc8051_siu_rtl.vhd:949:51  */
  assign n1558_o = s_recv_sh[7:1];
  assign n1559_o = {s_rxd_val, n1558_o};
  /* mc8051_siu_rtl.vhd:947:15  */
  assign n1560_o = s_m13_rxshift_en ? n1559_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:947:15  */
  assign n1563_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:946:13  */
  assign n1565_o = s_recv_state == 4'b0111;
  /* mc8051_siu_rtl.vhd:955:51  */
  assign n1566_o = s_recv_sh[7:1];
  assign n1567_o = {s_rxd_val, n1566_o};
  /* mc8051_siu_rtl.vhd:953:15  */
  assign n1568_o = s_m13_rxshift_en ? n1567_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:953:15  */
  assign n1571_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:952:13  */
  assign n1573_o = s_recv_state == 4'b1000;
  /* mc8051_siu_rtl.vhd:961:51  */
  assign n1574_o = s_recv_sh[7:1];
  assign n1575_o = {s_rxd_val, n1574_o};
  /* mc8051_siu_rtl.vhd:959:15  */
  assign n1576_o = s_m13_rxshift_en ? n1575_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:959:15  */
  assign n1579_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:958:13  */
  assign n1581_o = s_recv_state == 4'b1001;
  /* mc8051_siu_rtl.vhd:966:24  */
  assign n1582_o = ~s_ri;
  /* mc8051_siu_rtl.vhd:966:40  */
  assign n1583_o = ~s_sm2;
  /* mc8051_siu_rtl.vhd:966:30  */
  assign n1584_o = n1582_o & n1583_o;
  /* mc8051_siu_rtl.vhd:967:24  */
  assign n1585_o = ~s_ri;
  /* mc8051_siu_rtl.vhd:967:30  */
  assign n1586_o = n1585_o & s_rxd_val;
  /* mc8051_siu_rtl.vhd:966:47  */
  assign n1587_o = n1584_o | n1586_o;
  /* mc8051_siu_rtl.vhd:969:33  */
  assign n1588_o = s_rxpre_count[3:0];
  /* mc8051_siu_rtl.vhd:969:46  */
  assign n1590_o = n1588_o == 4'b1010;
  /* mc8051_siu_rtl.vhd:971:57  */
  assign n1591_o = s_recv_sh[7:1];
  /* mc8051_siu_rtl.vhd:966:15  */
  assign n1593_o = n1604_o ? 1'b1 : s_recv_done;
  /* mc8051_siu_rtl.vhd:966:15  */
  assign n1594_o = n1605_o ? s_rxd_val : s_rb8;
  assign n1595_o = {s_rxd_val, n1591_o};
  /* mc8051_siu_rtl.vhd:966:15  */
  assign n1596_o = n1606_o ? n1595_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:966:15  */
  assign n1597_o = n1607_o ? s_recv_sh : s_recv_buf;
  /* mc8051_siu_rtl.vhd:969:17  */
  assign n1600_o = n1590_o ? 2'b10 : 2'b00;
  /* mc8051_siu_rtl.vhd:979:17  */
  assign n1603_o = s_m13_rxshift_en ? 2'b10 : 2'b00;
  /* mc8051_siu_rtl.vhd:966:15  */
  assign n1604_o = n1587_o & n1590_o;
  /* mc8051_siu_rtl.vhd:966:15  */
  assign n1605_o = n1587_o & n1590_o;
  /* mc8051_siu_rtl.vhd:966:15  */
  assign n1606_o = n1587_o & n1590_o;
  /* mc8051_siu_rtl.vhd:966:15  */
  assign n1607_o = n1587_o & n1590_o;
  /* mc8051_siu_rtl.vhd:966:15  */
  assign n1608_o = n1587_o ? n1600_o : n1603_o;
  /* mc8051_siu_rtl.vhd:964:13  */
  assign n1610_o = s_recv_state == 4'b1010;
  assign n1611_o = {n1610_o, n1581_o, n1573_o, n1565_o, n1557_o, n1549_o, n1541_o, n1533_o, n1525_o, n1517_o, n1499_o};
  /* mc8051_siu_rtl.vhd:895:13  */
  always @*
    case (n1611_o)
      11'b10000000000: n1612_o = n1593_o;
      11'b01000000000: n1612_o = s_recv_done;
      11'b00100000000: n1612_o = s_recv_done;
      11'b00010000000: n1612_o = s_recv_done;
      11'b00001000000: n1612_o = s_recv_done;
      11'b00000100000: n1612_o = s_recv_done;
      11'b00000010000: n1612_o = s_recv_done;
      11'b00000001000: n1612_o = s_recv_done;
      11'b00000000100: n1612_o = s_recv_done;
      11'b00000000010: n1612_o = s_recv_done;
      11'b00000000001: n1612_o = n1492_o;
      default: n1612_o = s_recv_done;
    endcase
  /* mc8051_siu_rtl.vhd:895:13  */
  always @*
    case (n1611_o)
      11'b10000000000: n1613_o = n1594_o;
      11'b01000000000: n1613_o = s_rb8;
      11'b00100000000: n1613_o = s_rb8;
      11'b00010000000: n1613_o = s_rb8;
      11'b00001000000: n1613_o = s_rb8;
      11'b00000100000: n1613_o = s_rb8;
      11'b00000010000: n1613_o = s_rb8;
      11'b00000001000: n1613_o = s_rb8;
      11'b00000000100: n1613_o = s_rb8;
      11'b00000000010: n1613_o = s_rb8;
      11'b00000000001: n1613_o = s_rb8;
      default: n1613_o = s_rb8;
    endcase
  /* mc8051_siu_rtl.vhd:895:13  */
  always @*
    case (n1611_o)
      11'b10000000000: n1614_o = n1596_o;
      11'b01000000000: n1614_o = n1576_o;
      11'b00100000000: n1614_o = n1568_o;
      11'b00010000000: n1614_o = n1560_o;
      11'b00001000000: n1614_o = n1552_o;
      11'b00000100000: n1614_o = n1544_o;
      11'b00000010000: n1614_o = n1536_o;
      11'b00000001000: n1614_o = n1528_o;
      11'b00000000100: n1614_o = n1520_o;
      11'b00000000010: n1614_o = n1504_o;
      11'b00000000001: n1614_o = n1494_o;
      default: n1614_o = s_recv_sh;
    endcase
  /* mc8051_siu_rtl.vhd:895:13  */
  always @*
    case (n1611_o)
      11'b10000000000: n1615_o = n1597_o;
      11'b01000000000: n1615_o = s_recv_buf;
      11'b00100000000: n1615_o = s_recv_buf;
      11'b00010000000: n1615_o = s_recv_buf;
      11'b00001000000: n1615_o = s_recv_buf;
      11'b00000100000: n1615_o = s_recv_buf;
      11'b00000010000: n1615_o = s_recv_buf;
      11'b00000001000: n1615_o = s_recv_buf;
      11'b00000000100: n1615_o = s_recv_buf;
      11'b00000000010: n1615_o = s_recv_buf;
      11'b00000000001: n1615_o = s_recv_buf;
      default: n1615_o = s_recv_buf;
    endcase
  /* mc8051_siu_rtl.vhd:895:13  */
  always @*
    case (n1611_o)
      11'b10000000000: n1617_o = n1608_o;
      11'b01000000000: n1617_o = n1579_o;
      11'b00100000000: n1617_o = n1571_o;
      11'b00010000000: n1617_o = n1563_o;
      11'b00001000000: n1617_o = n1555_o;
      11'b00000100000: n1617_o = n1547_o;
      11'b00000010000: n1617_o = n1539_o;
      11'b00000001000: n1617_o = n1531_o;
      11'b00000000100: n1617_o = n1523_o;
      11'b00000000010: n1617_o = n1515_o;
      11'b00000000001: n1617_o = n1497_o;
      default: n1617_o = 2'b10;
    endcase
  /* mc8051_siu_rtl.vhd:894:11  */
  assign n1619_o = s_mode == 2'b01;
  /* mc8051_siu_rtl.vhd:993:30  */
  assign n1620_o = s_ren & s_detect;
  /* mc8051_siu_rtl.vhd:993:15  */
  assign n1622_o = n1620_o ? 1'b0 : s_recv_done;
  /* mc8051_siu_rtl.vhd:993:15  */
  assign n1624_o = n1620_o ? 8'b00000000 : s_recv_sh;
  /* mc8051_siu_rtl.vhd:993:15  */
  assign n1627_o = n1620_o ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:992:13  */
  assign n1629_o = s_recv_state == 4'b0000;
  /* mc8051_siu_rtl.vhd:999:28  */
  assign n1630_o = ~s_rxd_val;
  /* mc8051_siu_rtl.vhd:1002:53  */
  assign n1631_o = s_recv_sh[7:1];
  assign n1632_o = {s_rxd_val, n1631_o};
  /* mc8051_siu_rtl.vhd:999:15  */
  assign n1633_o = n1640_o ? n1632_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1000:17  */
  assign n1636_o = s_m2_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1006:17  */
  assign n1639_o = s_m2_rxshift_en ? 2'b10 : 2'b00;
  /* mc8051_siu_rtl.vhd:999:15  */
  assign n1640_o = n1630_o & s_m2_rxshift_en;
  /* mc8051_siu_rtl.vhd:999:15  */
  assign n1641_o = n1630_o ? n1636_o : n1639_o;
  /* mc8051_siu_rtl.vhd:998:13  */
  assign n1643_o = s_recv_state == 4'b0001;
  /* mc8051_siu_rtl.vhd:1013:51  */
  assign n1644_o = s_recv_sh[7:1];
  assign n1645_o = {s_rxd_val, n1644_o};
  /* mc8051_siu_rtl.vhd:1011:15  */
  assign n1646_o = s_m2_rxshift_en ? n1645_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1011:15  */
  assign n1649_o = s_m2_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1010:13  */
  assign n1651_o = s_recv_state == 4'b0010;
  /* mc8051_siu_rtl.vhd:1019:51  */
  assign n1652_o = s_recv_sh[7:1];
  assign n1653_o = {s_rxd_val, n1652_o};
  /* mc8051_siu_rtl.vhd:1017:15  */
  assign n1654_o = s_m2_rxshift_en ? n1653_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1017:15  */
  assign n1657_o = s_m2_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1016:13  */
  assign n1659_o = s_recv_state == 4'b0011;
  /* mc8051_siu_rtl.vhd:1025:51  */
  assign n1660_o = s_recv_sh[7:1];
  assign n1661_o = {s_rxd_val, n1660_o};
  /* mc8051_siu_rtl.vhd:1023:15  */
  assign n1662_o = s_m2_rxshift_en ? n1661_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1023:15  */
  assign n1665_o = s_m2_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1022:13  */
  assign n1667_o = s_recv_state == 4'b0100;
  /* mc8051_siu_rtl.vhd:1031:51  */
  assign n1668_o = s_recv_sh[7:1];
  assign n1669_o = {s_rxd_val, n1668_o};
  /* mc8051_siu_rtl.vhd:1029:15  */
  assign n1670_o = s_m2_rxshift_en ? n1669_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1029:15  */
  assign n1673_o = s_m2_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1028:13  */
  assign n1675_o = s_recv_state == 4'b0101;
  /* mc8051_siu_rtl.vhd:1037:51  */
  assign n1676_o = s_recv_sh[7:1];
  assign n1677_o = {s_rxd_val, n1676_o};
  /* mc8051_siu_rtl.vhd:1035:15  */
  assign n1678_o = s_m2_rxshift_en ? n1677_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1035:15  */
  assign n1681_o = s_m2_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1034:13  */
  assign n1683_o = s_recv_state == 4'b0110;
  /* mc8051_siu_rtl.vhd:1043:51  */
  assign n1684_o = s_recv_sh[7:1];
  assign n1685_o = {s_rxd_val, n1684_o};
  /* mc8051_siu_rtl.vhd:1041:15  */
  assign n1686_o = s_m2_rxshift_en ? n1685_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1041:15  */
  assign n1689_o = s_m2_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1040:13  */
  assign n1691_o = s_recv_state == 4'b0111;
  /* mc8051_siu_rtl.vhd:1049:51  */
  assign n1692_o = s_recv_sh[7:1];
  assign n1693_o = {s_rxd_val, n1692_o};
  /* mc8051_siu_rtl.vhd:1047:15  */
  assign n1694_o = s_m2_rxshift_en ? n1693_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1047:15  */
  assign n1697_o = s_m2_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1046:13  */
  assign n1699_o = s_recv_state == 4'b1000;
  /* mc8051_siu_rtl.vhd:1055:51  */
  assign n1700_o = s_recv_sh[7:1];
  assign n1701_o = {s_rxd_val, n1700_o};
  /* mc8051_siu_rtl.vhd:1053:15  */
  assign n1702_o = s_m2_rxshift_en ? n1701_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1053:15  */
  assign n1705_o = s_m2_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1052:13  */
  assign n1707_o = s_recv_state == 4'b1001;
  /* mc8051_siu_rtl.vhd:1060:24  */
  assign n1708_o = ~s_ri;
  /* mc8051_siu_rtl.vhd:1060:40  */
  assign n1709_o = ~s_sm2;
  /* mc8051_siu_rtl.vhd:1060:30  */
  assign n1710_o = n1708_o & n1709_o;
  /* mc8051_siu_rtl.vhd:1061:24  */
  assign n1711_o = ~s_ri;
  /* mc8051_siu_rtl.vhd:1061:30  */
  assign n1712_o = n1711_o & s_rxd_val;
  /* mc8051_siu_rtl.vhd:1060:47  */
  assign n1713_o = n1710_o | n1712_o;
  /* mc8051_siu_rtl.vhd:1064:53  */
  assign n1714_o = s_recv_sh[7:1];
  /* mc8051_siu_rtl.vhd:1060:15  */
  assign n1716_o = n1721_o ? 1'b1 : s_recv_done;
  /* mc8051_siu_rtl.vhd:1060:15  */
  assign n1717_o = n1722_o ? s_rxd_val : s_rb8;
  assign n1718_o = {s_rxd_val, n1714_o};
  /* mc8051_siu_rtl.vhd:1060:15  */
  assign n1719_o = n1723_o ? n1718_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1060:15  */
  assign n1720_o = n1724_o ? s_recv_sh : s_recv_buf;
  /* mc8051_siu_rtl.vhd:1060:15  */
  assign n1721_o = n1713_o & s_m2_rxshift_en;
  /* mc8051_siu_rtl.vhd:1060:15  */
  assign n1722_o = n1713_o & s_m2_rxshift_en;
  /* mc8051_siu_rtl.vhd:1060:15  */
  assign n1723_o = n1713_o & s_m2_rxshift_en;
  /* mc8051_siu_rtl.vhd:1060:15  */
  assign n1724_o = n1713_o & s_m2_rxshift_en;
  /* mc8051_siu_rtl.vhd:1071:15  */
  assign n1727_o = s_m2_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1058:13  */
  assign n1729_o = s_recv_state == 4'b1010;
  /* mc8051_siu_rtl.vhd:1076:15  */
  assign n1732_o = s_m2_rxshift_en ? 2'b10 : 2'b00;
  /* mc8051_siu_rtl.vhd:1074:13  */
  assign n1734_o = s_recv_state == 4'b1011;
  assign n1735_o = {n1734_o, n1729_o, n1707_o, n1699_o, n1691_o, n1683_o, n1675_o, n1667_o, n1659_o, n1651_o, n1643_o, n1629_o};
  /* mc8051_siu_rtl.vhd:991:13  */
  always @*
    case (n1735_o)
      12'b100000000000: n1736_o = s_recv_done;
      12'b010000000000: n1736_o = n1716_o;
      12'b001000000000: n1736_o = s_recv_done;
      12'b000100000000: n1736_o = s_recv_done;
      12'b000010000000: n1736_o = s_recv_done;
      12'b000001000000: n1736_o = s_recv_done;
      12'b000000100000: n1736_o = s_recv_done;
      12'b000000010000: n1736_o = s_recv_done;
      12'b000000001000: n1736_o = s_recv_done;
      12'b000000000100: n1736_o = s_recv_done;
      12'b000000000010: n1736_o = s_recv_done;
      12'b000000000001: n1736_o = n1622_o;
      default: n1736_o = s_recv_done;
    endcase
  /* mc8051_siu_rtl.vhd:991:13  */
  always @*
    case (n1735_o)
      12'b100000000000: n1737_o = s_rb8;
      12'b010000000000: n1737_o = n1717_o;
      12'b001000000000: n1737_o = s_rb8;
      12'b000100000000: n1737_o = s_rb8;
      12'b000010000000: n1737_o = s_rb8;
      12'b000001000000: n1737_o = s_rb8;
      12'b000000100000: n1737_o = s_rb8;
      12'b000000010000: n1737_o = s_rb8;
      12'b000000001000: n1737_o = s_rb8;
      12'b000000000100: n1737_o = s_rb8;
      12'b000000000010: n1737_o = s_rb8;
      12'b000000000001: n1737_o = s_rb8;
      default: n1737_o = s_rb8;
    endcase
  /* mc8051_siu_rtl.vhd:991:13  */
  always @*
    case (n1735_o)
      12'b100000000000: n1738_o = s_recv_sh;
      12'b010000000000: n1738_o = n1719_o;
      12'b001000000000: n1738_o = n1702_o;
      12'b000100000000: n1738_o = n1694_o;
      12'b000010000000: n1738_o = n1686_o;
      12'b000001000000: n1738_o = n1678_o;
      12'b000000100000: n1738_o = n1670_o;
      12'b000000010000: n1738_o = n1662_o;
      12'b000000001000: n1738_o = n1654_o;
      12'b000000000100: n1738_o = n1646_o;
      12'b000000000010: n1738_o = n1633_o;
      12'b000000000001: n1738_o = n1624_o;
      default: n1738_o = s_recv_sh;
    endcase
  /* mc8051_siu_rtl.vhd:991:13  */
  always @*
    case (n1735_o)
      12'b100000000000: n1739_o = s_recv_buf;
      12'b010000000000: n1739_o = n1720_o;
      12'b001000000000: n1739_o = s_recv_buf;
      12'b000100000000: n1739_o = s_recv_buf;
      12'b000010000000: n1739_o = s_recv_buf;
      12'b000001000000: n1739_o = s_recv_buf;
      12'b000000100000: n1739_o = s_recv_buf;
      12'b000000010000: n1739_o = s_recv_buf;
      12'b000000001000: n1739_o = s_recv_buf;
      12'b000000000100: n1739_o = s_recv_buf;
      12'b000000000010: n1739_o = s_recv_buf;
      12'b000000000001: n1739_o = s_recv_buf;
      default: n1739_o = s_recv_buf;
    endcase
  /* mc8051_siu_rtl.vhd:991:13  */
  always @*
    case (n1735_o)
      12'b100000000000: n1741_o = n1732_o;
      12'b010000000000: n1741_o = n1727_o;
      12'b001000000000: n1741_o = n1705_o;
      12'b000100000000: n1741_o = n1697_o;
      12'b000010000000: n1741_o = n1689_o;
      12'b000001000000: n1741_o = n1681_o;
      12'b000000100000: n1741_o = n1673_o;
      12'b000000010000: n1741_o = n1665_o;
      12'b000000001000: n1741_o = n1657_o;
      12'b000000000100: n1741_o = n1649_o;
      12'b000000000010: n1741_o = n1641_o;
      12'b000000000001: n1741_o = n1627_o;
      default: n1741_o = 2'b10;
    endcase
  /* mc8051_siu_rtl.vhd:990:11  */
  assign n1743_o = s_mode == 2'b10;
  /* mc8051_siu_rtl.vhd:1091:30  */
  assign n1744_o = s_ren & s_detect;
  /* mc8051_siu_rtl.vhd:1091:15  */
  assign n1746_o = n1744_o ? 1'b0 : s_recv_done;
  /* mc8051_siu_rtl.vhd:1091:15  */
  assign n1748_o = n1744_o ? 8'b00000000 : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1091:15  */
  assign n1751_o = n1744_o ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1090:13  */
  assign n1753_o = s_recv_state == 4'b0000;
  /* mc8051_siu_rtl.vhd:1097:27  */
  assign n1754_o = ~s_detect;
  /* mc8051_siu_rtl.vhd:1098:30  */
  assign n1755_o = ~s_rxd_val;
  /* mc8051_siu_rtl.vhd:1101:55  */
  assign n1756_o = s_recv_sh[7:1];
  assign n1757_o = {s_rxd_val, n1756_o};
  /* mc8051_siu_rtl.vhd:1097:15  */
  assign n1758_o = n1767_o ? n1757_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1099:19  */
  assign n1761_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1105:19  */
  assign n1764_o = s_m13_rxshift_en ? 2'b10 : 2'b00;
  /* mc8051_siu_rtl.vhd:1098:17  */
  assign n1765_o = n1755_o & s_m13_rxshift_en;
  /* mc8051_siu_rtl.vhd:1098:17  */
  assign n1766_o = n1755_o ? n1761_o : n1764_o;
  /* mc8051_siu_rtl.vhd:1097:15  */
  assign n1767_o = n1754_o & n1765_o;
  /* mc8051_siu_rtl.vhd:1097:15  */
  assign n1769_o = n1754_o ? n1766_o : 2'b00;
  /* mc8051_siu_rtl.vhd:1096:13  */
  assign n1771_o = s_recv_state == 4'b0001;
  /* mc8051_siu_rtl.vhd:1113:51  */
  assign n1772_o = s_recv_sh[7:1];
  assign n1773_o = {s_rxd_val, n1772_o};
  /* mc8051_siu_rtl.vhd:1111:15  */
  assign n1774_o = s_m13_rxshift_en ? n1773_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1111:15  */
  assign n1777_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1110:13  */
  assign n1779_o = s_recv_state == 4'b0010;
  /* mc8051_siu_rtl.vhd:1119:51  */
  assign n1780_o = s_recv_sh[7:1];
  assign n1781_o = {s_rxd_val, n1780_o};
  /* mc8051_siu_rtl.vhd:1117:15  */
  assign n1782_o = s_m13_rxshift_en ? n1781_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1117:15  */
  assign n1785_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1116:13  */
  assign n1787_o = s_recv_state == 4'b0011;
  /* mc8051_siu_rtl.vhd:1125:51  */
  assign n1788_o = s_recv_sh[7:1];
  assign n1789_o = {s_rxd_val, n1788_o};
  /* mc8051_siu_rtl.vhd:1123:15  */
  assign n1790_o = s_m13_rxshift_en ? n1789_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1123:15  */
  assign n1793_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1122:13  */
  assign n1795_o = s_recv_state == 4'b0100;
  /* mc8051_siu_rtl.vhd:1131:51  */
  assign n1796_o = s_recv_sh[7:1];
  assign n1797_o = {s_rxd_val, n1796_o};
  /* mc8051_siu_rtl.vhd:1129:15  */
  assign n1798_o = s_m13_rxshift_en ? n1797_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1129:15  */
  assign n1801_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1128:13  */
  assign n1803_o = s_recv_state == 4'b0101;
  /* mc8051_siu_rtl.vhd:1137:51  */
  assign n1804_o = s_recv_sh[7:1];
  assign n1805_o = {s_rxd_val, n1804_o};
  /* mc8051_siu_rtl.vhd:1135:15  */
  assign n1806_o = s_m13_rxshift_en ? n1805_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1135:15  */
  assign n1809_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1134:13  */
  assign n1811_o = s_recv_state == 4'b0110;
  /* mc8051_siu_rtl.vhd:1143:51  */
  assign n1812_o = s_recv_sh[7:1];
  assign n1813_o = {s_rxd_val, n1812_o};
  /* mc8051_siu_rtl.vhd:1141:15  */
  assign n1814_o = s_m13_rxshift_en ? n1813_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1141:15  */
  assign n1817_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1140:13  */
  assign n1819_o = s_recv_state == 4'b0111;
  /* mc8051_siu_rtl.vhd:1149:51  */
  assign n1820_o = s_recv_sh[7:1];
  assign n1821_o = {s_rxd_val, n1820_o};
  /* mc8051_siu_rtl.vhd:1147:15  */
  assign n1822_o = s_m13_rxshift_en ? n1821_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1147:15  */
  assign n1825_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1146:13  */
  assign n1827_o = s_recv_state == 4'b1000;
  /* mc8051_siu_rtl.vhd:1155:51  */
  assign n1828_o = s_recv_sh[7:1];
  assign n1829_o = {s_rxd_val, n1828_o};
  /* mc8051_siu_rtl.vhd:1153:15  */
  assign n1830_o = s_m13_rxshift_en ? n1829_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1153:15  */
  assign n1833_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1152:13  */
  assign n1835_o = s_recv_state == 4'b1001;
  /* mc8051_siu_rtl.vhd:1160:24  */
  assign n1836_o = ~s_ri;
  /* mc8051_siu_rtl.vhd:1160:40  */
  assign n1837_o = ~s_sm2;
  /* mc8051_siu_rtl.vhd:1160:30  */
  assign n1838_o = n1836_o & n1837_o;
  /* mc8051_siu_rtl.vhd:1161:24  */
  assign n1839_o = ~s_ri;
  /* mc8051_siu_rtl.vhd:1161:30  */
  assign n1840_o = n1839_o & s_rxd_val;
  /* mc8051_siu_rtl.vhd:1160:47  */
  assign n1841_o = n1838_o | n1840_o;
  /* mc8051_siu_rtl.vhd:1164:53  */
  assign n1842_o = s_recv_sh[7:1];
  /* mc8051_siu_rtl.vhd:1160:15  */
  assign n1844_o = n1849_o ? 1'b1 : s_recv_done;
  /* mc8051_siu_rtl.vhd:1160:15  */
  assign n1845_o = n1850_o ? s_rxd_val : s_rb8;
  assign n1846_o = {s_rxd_val, n1842_o};
  /* mc8051_siu_rtl.vhd:1160:15  */
  assign n1847_o = n1851_o ? n1846_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:1160:15  */
  assign n1848_o = n1852_o ? s_recv_sh : s_recv_buf;
  /* mc8051_siu_rtl.vhd:1160:15  */
  assign n1849_o = n1841_o & s_m13_rxshift_en;
  /* mc8051_siu_rtl.vhd:1160:15  */
  assign n1850_o = n1841_o & s_m13_rxshift_en;
  /* mc8051_siu_rtl.vhd:1160:15  */
  assign n1851_o = n1841_o & s_m13_rxshift_en;
  /* mc8051_siu_rtl.vhd:1160:15  */
  assign n1852_o = n1841_o & s_m13_rxshift_en;
  /* mc8051_siu_rtl.vhd:1171:15  */
  assign n1855_o = s_m13_rxshift_en ? 2'b01 : 2'b00;
  /* mc8051_siu_rtl.vhd:1158:13  */
  assign n1857_o = s_recv_state == 4'b1010;
  /* mc8051_siu_rtl.vhd:1176:15  */
  assign n1860_o = s_m13_rxshift_en ? 2'b10 : 2'b00;
  /* mc8051_siu_rtl.vhd:1174:13  */
  assign n1862_o = s_recv_state == 4'b1011;
  assign n1863_o = {n1862_o, n1857_o, n1835_o, n1827_o, n1819_o, n1811_o, n1803_o, n1795_o, n1787_o, n1779_o, n1771_o, n1753_o};
  /* mc8051_siu_rtl.vhd:1089:13  */
  always @*
    case (n1863_o)
      12'b100000000000: n1864_o = s_recv_done;
      12'b010000000000: n1864_o = n1844_o;
      12'b001000000000: n1864_o = s_recv_done;
      12'b000100000000: n1864_o = s_recv_done;
      12'b000010000000: n1864_o = s_recv_done;
      12'b000001000000: n1864_o = s_recv_done;
      12'b000000100000: n1864_o = s_recv_done;
      12'b000000010000: n1864_o = s_recv_done;
      12'b000000001000: n1864_o = s_recv_done;
      12'b000000000100: n1864_o = s_recv_done;
      12'b000000000010: n1864_o = s_recv_done;
      12'b000000000001: n1864_o = n1746_o;
      default: n1864_o = s_recv_done;
    endcase
  /* mc8051_siu_rtl.vhd:1089:13  */
  always @*
    case (n1863_o)
      12'b100000000000: n1865_o = s_rb8;
      12'b010000000000: n1865_o = n1845_o;
      12'b001000000000: n1865_o = s_rb8;
      12'b000100000000: n1865_o = s_rb8;
      12'b000010000000: n1865_o = s_rb8;
      12'b000001000000: n1865_o = s_rb8;
      12'b000000100000: n1865_o = s_rb8;
      12'b000000010000: n1865_o = s_rb8;
      12'b000000001000: n1865_o = s_rb8;
      12'b000000000100: n1865_o = s_rb8;
      12'b000000000010: n1865_o = s_rb8;
      12'b000000000001: n1865_o = s_rb8;
      default: n1865_o = s_rb8;
    endcase
  /* mc8051_siu_rtl.vhd:1089:13  */
  always @*
    case (n1863_o)
      12'b100000000000: n1866_o = s_recv_sh;
      12'b010000000000: n1866_o = n1847_o;
      12'b001000000000: n1866_o = n1830_o;
      12'b000100000000: n1866_o = n1822_o;
      12'b000010000000: n1866_o = n1814_o;
      12'b000001000000: n1866_o = n1806_o;
      12'b000000100000: n1866_o = n1798_o;
      12'b000000010000: n1866_o = n1790_o;
      12'b000000001000: n1866_o = n1782_o;
      12'b000000000100: n1866_o = n1774_o;
      12'b000000000010: n1866_o = n1758_o;
      12'b000000000001: n1866_o = n1748_o;
      default: n1866_o = s_recv_sh;
    endcase
  /* mc8051_siu_rtl.vhd:1089:13  */
  always @*
    case (n1863_o)
      12'b100000000000: n1867_o = s_recv_buf;
      12'b010000000000: n1867_o = n1848_o;
      12'b001000000000: n1867_o = s_recv_buf;
      12'b000100000000: n1867_o = s_recv_buf;
      12'b000010000000: n1867_o = s_recv_buf;
      12'b000001000000: n1867_o = s_recv_buf;
      12'b000000100000: n1867_o = s_recv_buf;
      12'b000000010000: n1867_o = s_recv_buf;
      12'b000000001000: n1867_o = s_recv_buf;
      12'b000000000100: n1867_o = s_recv_buf;
      12'b000000000010: n1867_o = s_recv_buf;
      12'b000000000001: n1867_o = s_recv_buf;
      default: n1867_o = s_recv_buf;
    endcase
  /* mc8051_siu_rtl.vhd:1089:13  */
  always @*
    case (n1863_o)
      12'b100000000000: n1869_o = n1860_o;
      12'b010000000000: n1869_o = n1855_o;
      12'b001000000000: n1869_o = n1833_o;
      12'b000100000000: n1869_o = n1825_o;
      12'b000010000000: n1869_o = n1817_o;
      12'b000001000000: n1869_o = n1809_o;
      12'b000000100000: n1869_o = n1801_o;
      12'b000000010000: n1869_o = n1793_o;
      12'b000000001000: n1869_o = n1785_o;
      12'b000000000100: n1869_o = n1777_o;
      12'b000000000010: n1869_o = n1769_o;
      12'b000000000001: n1869_o = n1751_o;
      default: n1869_o = 2'b10;
    endcase
  /* mc8051_siu_rtl.vhd:1088:11  */
  assign n1871_o = s_mode == 2'b11;
  assign n1872_o = {n1871_o, n1743_o, n1619_o, n1489_o};
  /* mc8051_siu_rtl.vhd:825:11  */
  always @*
    case (n1872_o)
      4'b1000: n1873_o = n1864_o;
      4'b0100: n1873_o = n1736_o;
      4'b0010: n1873_o = n1612_o;
      4'b0001: n1873_o = n1483_o;
      default: n1873_o = s_recv_done;
    endcase
  /* mc8051_siu_rtl.vhd:825:11  */
  always @*
    case (n1872_o)
      4'b1000: n1874_o = n1865_o;
      4'b0100: n1874_o = n1737_o;
      4'b0010: n1874_o = n1613_o;
      4'b0001: n1874_o = s_rb8;
      default: n1874_o = s_rb8;
    endcase
  /* mc8051_siu_rtl.vhd:825:11  */
  always @*
    case (n1872_o)
      4'b1000: n1875_o = n1866_o;
      4'b0100: n1875_o = n1738_o;
      4'b0010: n1875_o = n1614_o;
      4'b0001: n1875_o = n1484_o;
      default: n1875_o = s_recv_sh;
    endcase
  /* mc8051_siu_rtl.vhd:825:11  */
  always @*
    case (n1872_o)
      4'b1000: n1876_o = n1867_o;
      4'b0100: n1876_o = n1739_o;
      4'b0010: n1876_o = n1615_o;
      4'b0001: n1876_o = n1485_o;
      default: n1876_o = s_recv_buf;
    endcase
  /* mc8051_siu_rtl.vhd:825:11  */
  always @*
    case (n1872_o)
      4'b1000: n1878_o = n1869_o;
      4'b0100: n1878_o = n1741_o;
      4'b0010: n1878_o = n1617_o;
      4'b0001: n1878_o = n1487_o;
      default: n1878_o = 2'b00;
    endcase
  /* mc8051_siu_rtl.vhd:1188:44  */
  assign n1882_o = s_recv_state + 4'b0001;
  /* mc8051_siu_rtl.vhd:1187:13  */
  assign n1884_o = n1878_o == 2'b01;
  /* mc8051_siu_rtl.vhd:1189:13  */
  assign n1886_o = n1878_o == 2'b10;
  assign n1887_o = {n1886_o, n1884_o};
  /* mc8051_siu_rtl.vhd:1186:11  */
  always @*
    case (n1887_o)
      2'b10: n1889_o = 4'b0000;
      2'b01: n1889_o = n1882_o;
      default: n1889_o = s_recv_state;
    endcase
  /* mc8051_siu_rtl.vhd:213:9  */
  assign n1912_o = cen ? n604_o : s_rxpre_count;
  /* mc8051_siu_rtl.vhd:213:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1913_q <= 6'b000000;
    else
      n1913_q <= n1912_o;
  /* mc8051_siu_rtl.vhd:213:9  */
  assign n1914_o = cen ? n582_o : s_txpre_count;
  /* mc8051_siu_rtl.vhd:213:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1915_q <= 6'b000000;
    else
      n1915_q <= n1914_o;
  /* mc8051_siu_rtl.vhd:141:9  */
  assign n1916_o = cen ? tf_i : s_ff0;
  /* mc8051_siu_rtl.vhd:141:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1917_q <= 1'b0;
    else
      n1917_q <= n1916_o;
  /* mc8051_siu_rtl.vhd:141:9  */
  assign n1918_o = cen ? s_ff0 : s_ff1;
  /* mc8051_siu_rtl.vhd:141:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1919_q <= 1'b0;
    else
      n1919_q <= n1918_o;
  /* mc8051_siu_rtl.vhd:136:7  */
  assign n1920_o = {n475_o, n476_o};
  /* mc8051_siu_rtl.vhd:414:7  */
  assign n1921_o = cen ? n1356_o : s_txdm0;
  /* mc8051_siu_rtl.vhd:414:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1922_q <= 1'b1;
    else
      n1922_q <= n1921_o;
  /* mc8051_siu_rtl.vhd:141:9  */
  assign n1923_o = cen ? n506_o : s_trans;
  /* mc8051_siu_rtl.vhd:141:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1924_q <= 1'b0;
    else
      n1924_q <= n1923_o;
  /* mc8051_siu_rtl.vhd:819:9  */
  assign n1925_o = cen ? n1873_o : s_recv_done;
  /* mc8051_siu_rtl.vhd:819:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1926_q <= 1'b0;
    else
      n1926_q <= n1925_o;
  /* mc8051_siu_rtl.vhd:414:7  */
  assign n1927_o = cen ? n1357_o : s_tran_done;
  /* mc8051_siu_rtl.vhd:414:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1928_q <= 1'b0;
    else
      n1928_q <= n1927_o;
  /* mc8051_siu_rtl.vhd:819:9  */
  assign n1929_o = cen ? n1874_o : s_rb8;
  /* mc8051_siu_rtl.vhd:819:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1930_q <= 1'b0;
    else
      n1930_q <= n1929_o;
  /* mc8051_siu_rtl.vhd:819:9  */
  assign n1931_o = cen ? n1889_o : s_recv_state;
  /* mc8051_siu_rtl.vhd:819:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1932_q <= 4'b0000;
    else
      n1932_q <= n1931_o;
  /* mc8051_siu_rtl.vhd:414:7  */
  assign n1933_o = cen ? n1371_o : s_tran_state;
  /* mc8051_siu_rtl.vhd:414:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1934_q <= 4'b0000;
    else
      n1934_q <= n1933_o;
  /* mc8051_siu_rtl.vhd:305:7  */
  assign n1935_o = cen ? n770_o : s_rxd_ff0;
  /* mc8051_siu_rtl.vhd:305:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1936_q <= 1'b0;
    else
      n1936_q <= n1935_o;
  /* mc8051_siu_rtl.vhd:305:7  */
  assign n1937_o = cen ? n771_o : s_rxd_ff1;
  /* mc8051_siu_rtl.vhd:305:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1938_q <= 1'b0;
    else
      n1938_q <= n1937_o;
  /* mc8051_siu_rtl.vhd:305:7  */
  assign n1939_o = cen ? n772_o : s_rxd_ff2;
  /* mc8051_siu_rtl.vhd:305:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1940_q <= 1'b0;
    else
      n1940_q <= n1939_o;
  /* mc8051_siu_rtl.vhd:305:7  */
  assign n1941_o = cen ? n774_o : s_det_ff0;
  /* mc8051_siu_rtl.vhd:305:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1942_q <= 1'b0;
    else
      n1942_q <= n1941_o;
  /* mc8051_siu_rtl.vhd:305:7  */
  assign n1943_o = cen ? n776_o : s_det_ff1;
  /* mc8051_siu_rtl.vhd:305:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1944_q <= 1'b0;
    else
      n1944_q <= n1943_o;
  /* mc8051_siu_rtl.vhd:414:7  */
  assign n1945_o = cen ? n1358_o : s_tran_sh;
  /* mc8051_siu_rtl.vhd:414:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1946_q <= 11'b00000000000;
    else
      n1946_q <= n1945_o;
  /* mc8051_siu_rtl.vhd:819:9  */
  assign n1947_o = cen ? n1875_o : s_recv_sh;
  /* mc8051_siu_rtl.vhd:819:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1948_q <= 8'b00000000;
    else
      n1948_q <= n1947_o;
  /* mc8051_siu_rtl.vhd:819:9  */
  assign n1949_o = cen ? n1876_o : s_recv_buf;
  /* mc8051_siu_rtl.vhd:819:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1950_q <= 8'b00000000;
    else
      n1950_q <= n1949_o;
  /* mc8051_siu_rtl.vhd:213:9  */
  assign n1951_o = cen ? n617_o : s_rxm13_ff0;
  /* mc8051_siu_rtl.vhd:213:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1952_q <= 1'b0;
    else
      n1952_q <= n1951_o;
  /* mc8051_siu_rtl.vhd:213:9  */
  assign n1953_o = cen ? s_rxm13_ff0 : s_rxm13_ff1;
  /* mc8051_siu_rtl.vhd:213:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1954_q <= 1'b0;
    else
      n1954_q <= n1953_o;
  /* mc8051_siu_rtl.vhd:213:9  */
  assign n1955_o = cen ? n630_o : s_txm13_ff0;
  /* mc8051_siu_rtl.vhd:213:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1956_q <= 1'b0;
    else
      n1956_q <= n1955_o;
  /* mc8051_siu_rtl.vhd:213:9  */
  assign n1957_o = cen ? s_txm13_ff0 : s_txm13_ff1;
  /* mc8051_siu_rtl.vhd:213:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1958_q <= 1'b0;
    else
      n1958_q <= n1957_o;
  /* mc8051_siu_rtl.vhd:205:7  */
  assign n1959_o = {s_rb8, s_tran_done, s_recv_done};
  /* mc8051_siu_rtl.vhd:414:7  */
  assign n1960_o = cen ? n1351_o : n1961_q;
  /* mc8051_siu_rtl.vhd:414:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1961_q <= 1'b0;
    else
      n1961_q <= n1960_o;
  /* mc8051_siu_rtl.vhd:414:7  */
  assign n1962_o = cen ? n1355_o : n1963_q;
  /* mc8051_siu_rtl.vhd:414:7  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1963_q <= 1'b1;
    else
      n1963_q <= n1962_o;
endmodule

module mc8051_alu_8
  (input  [7:0] rom_data_i,
   input  [7:0] ram_data_i,
   input  [7:0] acc_i,
   input  [5:0] cmd_i,
   input  [1:0] cy_i,
   input  ov_i,
   output [1:0] new_cy_o,
   output new_ov_o,
   output [7:0] result_a_o,
   output [7:0] result_b_o);
  wire [7:0] s_alu_result;
  wire [1:0] s_alu_new_cy;
  wire [7:0] s_alu_op_a;
  wire [7:0] s_alu_op_b;
  wire [3:0] s_alu_cmd;
  wire [7:0] s_dvdnd;
  wire [7:0] s_dvsor;
  wire [7:0] s_qutnt;
  wire [7:0] s_rmndr;
  wire [7:0] s_mltplcnd;
  wire [7:0] s_mltplctr;
  wire [15:0] s_product;
  wire [7:0] s_dcml_data;
  wire [7:0] s_dcml_rslt;
  wire s_dcml_cy;
  wire [7:0] s_addsub_rslt;
  wire [1:0] s_addsub_newcy;
  wire s_addsub_ov;
  wire s_addsub_cy;
  wire s_addsub;
  wire [7:0] s_addsub_opa;
  wire [7:0] s_addsub_opb;
  wire [1:0] i_alumux_n392;
  wire i_alumux_n393;
  wire [7:0] i_alumux_n394;
  wire [7:0] i_alumux_n395;
  wire [7:0] i_alumux_n396;
  wire [7:0] i_alumux_n397;
  wire [3:0] i_alumux_n398;
  wire [7:0] i_alumux_n399;
  wire [7:0] i_alumux_n400;
  wire i_alumux_n401;
  wire i_alumux_n402;
  wire [7:0] i_alumux_n403;
  wire [7:0] i_alumux_n404;
  wire [7:0] i_alumux_n405;
  wire [7:0] i_alumux_n406;
  wire [7:0] i_alumux_n407;
  wire [1:0] i_alumux_cy_o;
  wire i_alumux_ov_o;
  wire [7:0] i_alumux_result_a_o;
  wire [7:0] i_alumux_result_b_o;
  wire [7:0] i_alumux_op_a_o;
  wire [7:0] i_alumux_op_b_o;
  wire [3:0] i_alumux_alu_cmd_o;
  wire [7:0] i_alumux_opa_o;
  wire [7:0] i_alumux_opb_o;
  wire i_alumux_addsub_o;
  wire i_alumux_addsub_cy_o;
  wire [7:0] i_alumux_dvdnd_o;
  wire [7:0] i_alumux_dvsor_o;
  wire [7:0] i_alumux_mltplcnd_o;
  wire [7:0] i_alumux_mltplctr_o;
  wire [7:0] i_alumux_dcml_data_o;
  wire [1:0] i_alucore_n440;
  wire [7:0] i_alucore_n441;
  wire [1:0] i_alucore_cy_o;
  wire [7:0] i_alucore_result_o;
  wire [1:0] i_addsub_core_n446;
  wire i_addsub_core_n447;
  wire [7:0] i_addsub_core_n448;
  wire [1:0] i_addsub_core_cy_o;
  wire i_addsub_core_ov_o;
  wire [7:0] i_addsub_core_rslt_o;
  wire [15:0] gen_multiplier1_i_comb_mltplr_n455;
  wire [15:0] gen_multiplier1_i_comb_mltplr_product_o;
  wire [7:0] gen_divider1_i_comb_divider_n458;
  wire [7:0] gen_divider1_i_comb_divider_n459;
  wire [7:0] gen_divider1_i_comb_divider_qutnt_o;
  wire [7:0] gen_divider1_i_comb_divider_rmndr_o;
  wire [7:0] gen_dcml_adj1_i_dcml_adjust_n464;
  wire gen_dcml_adj1_i_dcml_adjust_n465;
  wire [7:0] gen_dcml_adj1_i_dcml_adjust_data_o;
  wire gen_dcml_adj1_i_dcml_adjust_cy_o;
  assign new_cy_o = i_alumux_n392;
  assign new_ov_o = i_alumux_n393;
  assign result_a_o = i_alumux_n394;
  assign result_b_o = i_alumux_n395;
  /* mc8051_alu_struc.vhd:69:10  */
  assign s_alu_result = i_alucore_n441; // (signal)
  /* mc8051_alu_struc.vhd:70:10  */
  assign s_alu_new_cy = i_alucore_n440; // (signal)
  /* mc8051_alu_struc.vhd:71:10  */
  assign s_alu_op_a = i_alumux_n396; // (signal)
  /* mc8051_alu_struc.vhd:72:10  */
  assign s_alu_op_b = i_alumux_n397; // (signal)
  /* mc8051_alu_struc.vhd:73:10  */
  assign s_alu_cmd = i_alumux_n398; // (signal)
  /* mc8051_alu_struc.vhd:74:10  */
  assign s_dvdnd = i_alumux_n403; // (signal)
  /* mc8051_alu_struc.vhd:75:10  */
  assign s_dvsor = i_alumux_n404; // (signal)
  /* mc8051_alu_struc.vhd:76:10  */
  assign s_qutnt = gen_divider1_i_comb_divider_n458; // (signal)
  /* mc8051_alu_struc.vhd:77:10  */
  assign s_rmndr = gen_divider1_i_comb_divider_n459; // (signal)
  /* mc8051_alu_struc.vhd:78:10  */
  assign s_mltplcnd = i_alumux_n405; // (signal)
  /* mc8051_alu_struc.vhd:79:10  */
  assign s_mltplctr = i_alumux_n406; // (signal)
  /* mc8051_alu_struc.vhd:80:10  */
  assign s_product = gen_multiplier1_i_comb_mltplr_n455; // (signal)
  /* mc8051_alu_struc.vhd:81:10  */
  assign s_dcml_data = i_alumux_n407; // (signal)
  /* mc8051_alu_struc.vhd:82:10  */
  assign s_dcml_rslt = gen_dcml_adj1_i_dcml_adjust_n464; // (signal)
  /* mc8051_alu_struc.vhd:83:10  */
  assign s_dcml_cy = gen_dcml_adj1_i_dcml_adjust_n465; // (signal)
  /* mc8051_alu_struc.vhd:84:10  */
  assign s_addsub_rslt = i_addsub_core_n448; // (signal)
  /* mc8051_alu_struc.vhd:85:10  */
  assign s_addsub_newcy = i_addsub_core_n446; // (signal)
  /* mc8051_alu_struc.vhd:86:10  */
  assign s_addsub_ov = i_addsub_core_n447; // (signal)
  /* mc8051_alu_struc.vhd:87:10  */
  assign s_addsub_cy = i_alumux_n402; // (signal)
  /* mc8051_alu_struc.vhd:88:10  */
  assign s_addsub = i_alumux_n401; // (signal)
  /* mc8051_alu_struc.vhd:89:10  */
  assign s_addsub_opa = i_alumux_n399; // (signal)
  /* mc8051_alu_struc.vhd:90:10  */
  assign s_addsub_opb = i_alumux_n400; // (signal)
  /* mc8051_alu_struc.vhd:105:24  */
  assign i_alumux_n392 = i_alumux_cy_o; // (signal)
  /* mc8051_alu_struc.vhd:106:24  */
  assign i_alumux_n393 = i_alumux_ov_o; // (signal)
  /* mc8051_alu_struc.vhd:107:24  */
  assign i_alumux_n394 = i_alumux_result_a_o; // (signal)
  /* mc8051_alu_struc.vhd:108:24  */
  assign i_alumux_n395 = i_alumux_result_b_o; // (signal)
  /* mc8051_alu_struc.vhd:115:24  */
  assign i_alumux_n396 = i_alumux_op_a_o; // (signal)
  /* mc8051_alu_struc.vhd:116:24  */
  assign i_alumux_n397 = i_alumux_op_b_o; // (signal)
  /* mc8051_alu_struc.vhd:117:24  */
  assign i_alumux_n398 = i_alumux_alu_cmd_o; // (signal)
  /* mc8051_alu_struc.vhd:118:24  */
  assign i_alumux_n399 = i_alumux_opa_o; // (signal)
  /* mc8051_alu_struc.vhd:119:24  */
  assign i_alumux_n400 = i_alumux_opb_o; // (signal)
  /* mc8051_alu_struc.vhd:120:24  */
  assign i_alumux_n401 = i_alumux_addsub_o; // (signal)
  /* mc8051_alu_struc.vhd:121:24  */
  assign i_alumux_n402 = i_alumux_addsub_cy_o; // (signal)
  /* mc8051_alu_struc.vhd:122:24  */
  assign i_alumux_n403 = i_alumux_dvdnd_o; // (signal)
  /* mc8051_alu_struc.vhd:123:24  */
  assign i_alumux_n404 = i_alumux_dvsor_o; // (signal)
  /* mc8051_alu_struc.vhd:126:24  */
  assign i_alumux_n405 = i_alumux_mltplcnd_o; // (signal)
  /* mc8051_alu_struc.vhd:127:24  */
  assign i_alumux_n406 = i_alumux_mltplctr_o; // (signal)
  /* mc8051_alu_struc.vhd:129:24  */
  assign i_alumux_n407 = i_alumux_dcml_data_o; // (signal)
  /* mc8051_alu_struc.vhd:94:3  */
  alumux_8 i_alumux (
    .rom_data_i(rom_data_i),
    .ram_data_i(ram_data_i),
    .acc_i(acc_i),
    .cmd_i(cmd_i),
    .cy_i(cy_i),
    .ov_i(ov_i),
    .result_i(s_alu_result),
    .new_cy_i(s_alu_new_cy),
    .addsub_rslt_i(s_addsub_rslt),
    .addsub_cy_i(s_addsub_newcy),
    .addsub_ov_i(s_addsub_ov),
    .qutnt_i(s_qutnt),
    .rmndr_i(s_rmndr),
    .product_i(s_product),
    .dcml_data_i(s_dcml_rslt),
    .dcml_cy_i(s_dcml_cy),
    .cy_o(i_alumux_cy_o),
    .ov_o(i_alumux_ov_o),
    .result_a_o(i_alumux_result_a_o),
    .result_b_o(i_alumux_result_b_o),
    .op_a_o(i_alumux_op_a_o),
    .op_b_o(i_alumux_op_b_o),
    .alu_cmd_o(i_alumux_alu_cmd_o),
    .opa_o(i_alumux_opa_o),
    .opb_o(i_alumux_opb_o),
    .addsub_o(i_alumux_addsub_o),
    .addsub_cy_o(i_alumux_addsub_cy_o),
    .dvdnd_o(i_alumux_dvdnd_o),
    .dvsor_o(i_alumux_dvsor_o),
    .mltplcnd_o(i_alumux_mltplcnd_o),
    .mltplctr_o(i_alumux_mltplctr_o),
    .dcml_data_o(i_alumux_dcml_data_o));
  /* mc8051_alu_struc.vhd:141:20  */
  assign i_alucore_n440 = i_alucore_cy_o; // (signal)
  /* mc8051_alu_struc.vhd:142:20  */
  assign i_alucore_n441 = i_alucore_result_o; // (signal)
  /* mc8051_alu_struc.vhd:133:3  */
  alucore_8 i_alucore (
    .op_a_i(s_alu_op_a),
    .op_b_i(s_alu_op_b),
    .alu_cmd_i(s_alu_cmd),
    .cy_i(cy_i),
    .cy_o(i_alucore_cy_o),
    .result_o(i_alucore_result_o));
  /* mc8051_alu_struc.vhd:150:27  */
  assign i_addsub_core_n446 = i_addsub_core_cy_o; // (signal)
  /* mc8051_alu_struc.vhd:151:27  */
  assign i_addsub_core_n447 = i_addsub_core_ov_o; // (signal)
  /* mc8051_alu_struc.vhd:152:27  */
  assign i_addsub_core_n448 = i_addsub_core_rslt_o; // (signal)
  /* mc8051_alu_struc.vhd:144:3  */
  addsub_core_8 i_addsub_core (
    .opa_i(s_addsub_opa),
    .opb_i(s_addsub_opb),
    .addsub_i(s_addsub),
    .cy_i(s_addsub_cy),
    .cy_o(i_addsub_core_cy_o),
    .ov_o(i_addsub_core_ov_o),
    .rslt_o(i_addsub_core_rslt_o));
  /* mc8051_alu_struc.vhd:161:23  */
  assign gen_multiplier1_i_comb_mltplr_n455 = gen_multiplier1_i_comb_mltplr_product_o; // (signal)
  /* mc8051_alu_struc.vhd:155:5  */
  comb_mltplr_8 gen_multiplier1_i_comb_mltplr (
    .mltplcnd_i(s_mltplcnd),
    .mltplctr_i(s_mltplctr),
    .product_o(gen_multiplier1_i_comb_mltplr_product_o));
  /* mc8051_alu_struc.vhd:174:20  */
  assign gen_divider1_i_comb_divider_n458 = gen_divider1_i_comb_divider_qutnt_o; // (signal)
  /* mc8051_alu_struc.vhd:175:20  */
  assign gen_divider1_i_comb_divider_n459 = gen_divider1_i_comb_divider_rmndr_o; // (signal)
  /* mc8051_alu_struc.vhd:168:5  */
  comb_divider_8 gen_divider1_i_comb_divider (
    .dvdnd_i(s_dvdnd),
    .dvsor_i(s_dvsor),
    .qutnt_o(gen_divider1_i_comb_divider_qutnt_o),
    .rmndr_o(gen_divider1_i_comb_divider_rmndr_o));
  /* mc8051_alu_struc.vhd:189:19  */
  assign gen_dcml_adj1_i_dcml_adjust_n464 = gen_dcml_adj1_i_dcml_adjust_data_o; // (signal)
  /* mc8051_alu_struc.vhd:190:19  */
  assign gen_dcml_adj1_i_dcml_adjust_n465 = gen_dcml_adj1_i_dcml_adjust_cy_o; // (signal)
  /* mc8051_alu_struc.vhd:183:5  */
  dcml_adjust_8 gen_dcml_adj1_i_dcml_adjust (
    .data_i(s_dcml_data),
    .cy_i(cy_i),
    .data_o(gen_dcml_adj1_i_dcml_adjust_data_o),
    .cy_o(gen_dcml_adj1_i_dcml_adjust_cy_o));
endmodule

module mc8051_control
  (input  [7:0] rom_data_i,
   input  [7:0] ram_data_i,
   input  [7:0] aludata_i,
   input  [7:0] aludatb_i,
   input  [1:0] new_cy_i,
   input  new_ov_i,
   input  reset,
   input  clk,
   input  cen,
   input  int0_i,
   input  int1_i,
   input  [7:0] datax_i,
   input  [7:0] p0_i,
   input  [7:0] p1_i,
   input  [7:0] p2_i,
   input  [7:0] p3_i,
   input  [2:0] all_scon_i,
   input  [7:0] all_sbuf_i,
   input  all_tf0_i,
   input  all_tf1_i,
   input  [7:0] all_tl0_i,
   input  [7:0] all_tl1_i,
   input  [7:0] all_th0_i,
   input  [7:0] all_th1_i,
   output [15:0] pc_o,
   output [7:0] ram_data_o,
   output [6:0] ram_adr_o,
   output [7:0] reg_data_o,
   output ram_wr_o,
   output [1:0] cy_o,
   output ov_o,
   output ram_en_o,
   output [5:0] alu_cmd_o,
   output [7:0] acc_o,
   output [7:0] datax_o,
   output [15:0] adrx_o,
   output wrx_o,
   output memx_o,
   output [7:0] p0_o,
   output [7:0] p1_o,
   output [7:0] p2_o,
   output [7:0] p3_o,
   output all_trans_o,
   output [5:0] all_scon_o,
   output [7:0] all_sbuf_o,
   output all_smod_o,
   output all_tcon_tr0_o,
   output all_tcon_tr1_o,
   output [7:0] all_tmod_o,
   output [7:0] all_reload_o,
   output [1:0] all_wt_o,
   output all_wt_en_o);
  wire [3:0] s_pc_inc_en;
  wire [2:0] s_regs_wr_en;
  wire [3:0] s_data_mux;
  wire [3:0] s_bdata_mux;
  wire [3:0] s_adr_mux;
  wire [1:0] s_adrx_mux;
  wire s_wrx_mux;
  wire [3:0] s_help_en;
  wire [1:0] s_help16_en;
  wire s_helpb_en;
  wire s_intpre2_d;
  wire s_intpre2_en;
  wire s_intlow_d;
  wire s_intlow_en;
  wire s_inthigh_d;
  wire s_inthigh_en;
  wire [2:0] s_nextstate;
  wire [2:0] state;
  wire [7:0] s_command;
  wire [7:0] s_help;
  wire s_bit_data;
  wire s_intpre;
  wire s_intpre2;
  wire s_inthigh;
  wire s_intlow;
  wire s_intblock;
  wire s_ri;
  wire s_ti;
  wire s_tf1;
  wire s_tf0;
  wire s_ie1;
  wire s_ie0;
  wire [7:0] ie;
  wire [7:0] ip;
  wire [7:0] psw;
  wire [7:0] acc;
  wire s_ext0isr_d;
  wire s_ext1isr_d;
  wire s_ext0isrh_d;
  wire s_ext1isrh_d;
  wire s_ext0isr_en;
  wire s_ext1isr_en;
  wire s_ext0isrh_en;
  wire s_ext1isrh_en;
  wire [5:0] i_control_fsm_n175;
  wire [3:0] i_control_fsm_n176;
  wire [2:0] i_control_fsm_n177;
  wire [3:0] i_control_fsm_n178;
  wire [1:0] i_control_fsm_n179;
  wire i_control_fsm_n180;
  wire [3:0] i_control_fsm_n181;
  wire [3:0] i_control_fsm_n182;
  wire [2:0] i_control_fsm_n183;
  wire [3:0] i_control_fsm_n184;
  wire [1:0] i_control_fsm_n185;
  wire i_control_fsm_n186;
  wire i_control_fsm_n187;
  wire i_control_fsm_n188;
  wire i_control_fsm_n189;
  wire i_control_fsm_n190;
  wire i_control_fsm_n191;
  wire i_control_fsm_n192;
  wire i_control_fsm_n193;
  wire i_control_fsm_n194;
  wire i_control_fsm_n195;
  wire i_control_fsm_n196;
  wire i_control_fsm_n197;
  wire i_control_fsm_n198;
  wire i_control_fsm_n199;
  wire i_control_fsm_n200;
  wire [5:0] i_control_fsm_alu_cmd_o;
  wire [3:0] i_control_fsm_pc_inc_en_o;
  wire [2:0] i_control_fsm_nextstate_o;
  wire [3:0] i_control_fsm_adr_mux_o;
  wire [1:0] i_control_fsm_adrx_mux_o;
  wire i_control_fsm_wrx_mux_o;
  wire [3:0] i_control_fsm_data_mux_o;
  wire [3:0] i_control_fsm_bdata_mux_o;
  wire [2:0] i_control_fsm_regs_wr_en_o;
  wire [3:0] i_control_fsm_help_en_o;
  wire [1:0] i_control_fsm_help16_en_o;
  wire i_control_fsm_helpb_en_o;
  wire i_control_fsm_inthigh_en_o;
  wire i_control_fsm_intlow_en_o;
  wire i_control_fsm_intpre2_en_o;
  wire i_control_fsm_inthigh_d_o;
  wire i_control_fsm_intlow_d_o;
  wire i_control_fsm_intpre2_d_o;
  wire i_control_fsm_ext0isr_d_o;
  wire i_control_fsm_ext1isr_d_o;
  wire i_control_fsm_ext0isrh_d_o;
  wire i_control_fsm_ext1isrh_d_o;
  wire i_control_fsm_ext0isr_en_o;
  wire i_control_fsm_ext1isr_en_o;
  wire i_control_fsm_ext0isrh_en_o;
  wire i_control_fsm_ext1isrh_en_o;
  wire [15:0] i_control_mem_n253;
  wire [7:0] i_control_mem_n254;
  wire [6:0] i_control_mem_n255;
  wire [7:0] i_control_mem_n256;
  wire i_control_mem_n257;
  wire [1:0] i_control_mem_n258;
  wire i_control_mem_n259;
  wire i_control_mem_n260;
  wire [7:0] i_control_mem_n261;
  wire [7:0] i_control_mem_n262;
  wire [7:0] i_control_mem_n263;
  wire [7:0] i_control_mem_n264;
  wire [7:0] i_control_mem_n265;
  wire i_control_mem_n266;
  wire [5:0] i_control_mem_n267;
  wire [7:0] i_control_mem_n268;
  wire i_control_mem_n269;
  wire i_control_mem_n270;
  wire i_control_mem_n271;
  wire [7:0] i_control_mem_n272;
  wire [7:0] i_control_mem_n273;
  wire [1:0] i_control_mem_n274;
  wire i_control_mem_n275;
  wire [2:0] i_control_mem_n276;
  wire [7:0] i_control_mem_n277;
  wire i_control_mem_n278;
  wire [7:0] i_control_mem_n279;
  wire i_control_mem_n280;
  wire i_control_mem_n281;
  wire i_control_mem_n282;
  wire i_control_mem_n283;
  wire i_control_mem_n284;
  wire i_control_mem_n285;
  wire i_control_mem_n286;
  wire i_control_mem_n287;
  wire i_control_mem_n288;
  wire i_control_mem_n289;
  wire i_control_mem_n290;
  wire [7:0] i_control_mem_n291;
  wire [7:0] i_control_mem_n292;
  wire [7:0] i_control_mem_n293;
  wire [15:0] i_control_mem_n294;
  wire [7:0] i_control_mem_n295;
  wire i_control_mem_n296;
  wire i_control_mem_n297;
  wire [15:0] i_control_mem_pc_o;
  wire [7:0] i_control_mem_ram_data_o;
  wire [6:0] i_control_mem_ram_adr_o;
  wire [7:0] i_control_mem_reg_data_o;
  wire i_control_mem_ram_wr_o;
  wire [1:0] i_control_mem_cy_o;
  wire i_control_mem_ov_o;
  wire i_control_mem_ram_en_o;
  wire [7:0] i_control_mem_acc_o;
  wire [7:0] i_control_mem_p0_o;
  wire [7:0] i_control_mem_p1_o;
  wire [7:0] i_control_mem_p2_o;
  wire [7:0] i_control_mem_p3_o;
  wire i_control_mem_all_trans_o;
  wire [5:0] i_control_mem_all_scon_o;
  wire [7:0] i_control_mem_all_sbuf_o;
  wire i_control_mem_all_smod_o;
  wire i_control_mem_all_tcon_tr0_o;
  wire i_control_mem_all_tcon_tr1_o;
  wire [7:0] i_control_mem_all_tmod_o;
  wire [7:0] i_control_mem_all_reload_o;
  wire [1:0] i_control_mem_all_wt_o;
  wire i_control_mem_all_wt_en_o;
  wire [2:0] i_control_mem_state_o;
  wire [7:0] i_control_mem_help_o;
  wire i_control_mem_bit_data_o;
  wire [7:0] i_control_mem_command_o;
  wire i_control_mem_inthigh_o;
  wire i_control_mem_intlow_o;
  wire i_control_mem_intpre_o;
  wire i_control_mem_intpre2_o;
  wire i_control_mem_intblock_o;
  wire i_control_mem_ti_o;
  wire i_control_mem_ri_o;
  wire i_control_mem_ie0_o;
  wire i_control_mem_ie1_o;
  wire i_control_mem_tf0_o;
  wire i_control_mem_tf1_o;
  wire [7:0] i_control_mem_psw_o;
  wire [7:0] i_control_mem_ie_o;
  wire [7:0] i_control_mem_ip_o;
  wire [15:0] i_control_mem_adrx_o;
  wire [7:0] i_control_mem_datax_o;
  wire i_control_mem_wrx_o;
  wire i_control_mem_memx_o;
  assign pc_o = i_control_mem_n253;
  assign ram_data_o = i_control_mem_n254;
  assign ram_adr_o = i_control_mem_n255;
  assign reg_data_o = i_control_mem_n256;
  assign ram_wr_o = i_control_mem_n257;
  assign cy_o = i_control_mem_n258;
  assign ov_o = i_control_mem_n259;
  assign ram_en_o = i_control_mem_n260;
  assign alu_cmd_o = i_control_fsm_n175;
  assign acc_o = acc;
  assign datax_o = i_control_mem_n295;
  assign adrx_o = i_control_mem_n294;
  assign wrx_o = i_control_mem_n297;
  assign memx_o = i_control_mem_n296;
  assign p0_o = i_control_mem_n262;
  assign p1_o = i_control_mem_n263;
  assign p2_o = i_control_mem_n264;
  assign p3_o = i_control_mem_n265;
  assign all_trans_o = i_control_mem_n266;
  assign all_scon_o = i_control_mem_n267;
  assign all_sbuf_o = i_control_mem_n268;
  assign all_smod_o = i_control_mem_n269;
  assign all_tcon_tr0_o = i_control_mem_n270;
  assign all_tcon_tr1_o = i_control_mem_n271;
  assign all_tmod_o = i_control_mem_n272;
  assign all_reload_o = i_control_mem_n273;
  assign all_wt_o = i_control_mem_n274;
  assign all_wt_en_o = i_control_mem_n275;
  /* mc8051_control_struc.vhd:70:10  */
  assign s_pc_inc_en = i_control_fsm_n176; // (signal)
  /* mc8051_control_struc.vhd:71:10  */
  assign s_regs_wr_en = i_control_fsm_n183; // (signal)
  /* mc8051_control_struc.vhd:72:10  */
  assign s_data_mux = i_control_fsm_n181; // (signal)
  /* mc8051_control_struc.vhd:73:10  */
  assign s_bdata_mux = i_control_fsm_n182; // (signal)
  /* mc8051_control_struc.vhd:74:10  */
  assign s_adr_mux = i_control_fsm_n178; // (signal)
  /* mc8051_control_struc.vhd:75:10  */
  assign s_adrx_mux = i_control_fsm_n179; // (signal)
  /* mc8051_control_struc.vhd:76:10  */
  assign s_wrx_mux = i_control_fsm_n180; // (signal)
  /* mc8051_control_struc.vhd:77:10  */
  assign s_help_en = i_control_fsm_n184; // (signal)
  /* mc8051_control_struc.vhd:78:10  */
  assign s_help16_en = i_control_fsm_n185; // (signal)
  /* mc8051_control_struc.vhd:79:10  */
  assign s_helpb_en = i_control_fsm_n186; // (signal)
  /* mc8051_control_struc.vhd:80:10  */
  assign s_intpre2_d = i_control_fsm_n192; // (signal)
  /* mc8051_control_struc.vhd:81:10  */
  assign s_intpre2_en = i_control_fsm_n189; // (signal)
  /* mc8051_control_struc.vhd:82:10  */
  assign s_intlow_d = i_control_fsm_n191; // (signal)
  /* mc8051_control_struc.vhd:83:10  */
  assign s_intlow_en = i_control_fsm_n188; // (signal)
  /* mc8051_control_struc.vhd:84:10  */
  assign s_inthigh_d = i_control_fsm_n190; // (signal)
  /* mc8051_control_struc.vhd:85:10  */
  assign s_inthigh_en = i_control_fsm_n187; // (signal)
  /* mc8051_control_struc.vhd:86:10  */
  assign s_nextstate = i_control_fsm_n177; // (signal)
  /* mc8051_control_struc.vhd:87:10  */
  assign state = i_control_mem_n276; // (signal)
  /* mc8051_control_struc.vhd:88:10  */
  assign s_command = i_control_mem_n279; // (signal)
  /* mc8051_control_struc.vhd:89:10  */
  assign s_help = i_control_mem_n277; // (signal)
  /* mc8051_control_struc.vhd:90:10  */
  assign s_bit_data = i_control_mem_n278; // (signal)
  /* mc8051_control_struc.vhd:91:10  */
  assign s_intpre = i_control_mem_n282; // (signal)
  /* mc8051_control_struc.vhd:92:10  */
  assign s_intpre2 = i_control_mem_n283; // (signal)
  /* mc8051_control_struc.vhd:93:10  */
  assign s_inthigh = i_control_mem_n280; // (signal)
  /* mc8051_control_struc.vhd:94:10  */
  assign s_intlow = i_control_mem_n281; // (signal)
  /* mc8051_control_struc.vhd:95:10  */
  assign s_intblock = i_control_mem_n284; // (signal)
  /* mc8051_control_struc.vhd:96:10  */
  assign s_ri = i_control_mem_n286; // (signal)
  /* mc8051_control_struc.vhd:97:10  */
  assign s_ti = i_control_mem_n285; // (signal)
  /* mc8051_control_struc.vhd:98:10  */
  assign s_tf1 = i_control_mem_n290; // (signal)
  /* mc8051_control_struc.vhd:99:10  */
  assign s_tf0 = i_control_mem_n289; // (signal)
  /* mc8051_control_struc.vhd:100:10  */
  assign s_ie1 = i_control_mem_n288; // (signal)
  /* mc8051_control_struc.vhd:101:10  */
  assign s_ie0 = i_control_mem_n287; // (signal)
  /* mc8051_control_struc.vhd:102:10  */
  assign ie = i_control_mem_n292; // (signal)
  /* mc8051_control_struc.vhd:103:10  */
  assign ip = i_control_mem_n293; // (signal)
  /* mc8051_control_struc.vhd:104:10  */
  assign psw = i_control_mem_n291; // (signal)
  /* mc8051_control_struc.vhd:105:10  */
  assign acc = i_control_mem_n261; // (signal)
  /* mc8051_control_struc.vhd:106:10  */
  assign s_ext0isr_d = i_control_fsm_n193; // (signal)
  /* mc8051_control_struc.vhd:107:10  */
  assign s_ext1isr_d = i_control_fsm_n194; // (signal)
  /* mc8051_control_struc.vhd:108:10  */
  assign s_ext0isrh_d = i_control_fsm_n195; // (signal)
  /* mc8051_control_struc.vhd:109:10  */
  assign s_ext1isrh_d = i_control_fsm_n196; // (signal)
  /* mc8051_control_struc.vhd:110:10  */
  assign s_ext0isr_en = i_control_fsm_n197; // (signal)
  /* mc8051_control_struc.vhd:111:10  */
  assign s_ext1isr_en = i_control_fsm_n198; // (signal)
  /* mc8051_control_struc.vhd:112:10  */
  assign s_ext0isrh_en = i_control_fsm_n199; // (signal)
  /* mc8051_control_struc.vhd:113:10  */
  assign s_ext1isrh_en = i_control_fsm_n200; // (signal)
  /* mc8051_control_struc.vhd:143:30  */
  assign i_control_fsm_n175 = i_control_fsm_alu_cmd_o; // (signal)
  /* mc8051_control_struc.vhd:144:30  */
  assign i_control_fsm_n176 = i_control_fsm_pc_inc_en_o; // (signal)
  /* mc8051_control_struc.vhd:145:30  */
  assign i_control_fsm_n177 = i_control_fsm_nextstate_o; // (signal)
  /* mc8051_control_struc.vhd:146:30  */
  assign i_control_fsm_n178 = i_control_fsm_adr_mux_o; // (signal)
  /* mc8051_control_struc.vhd:147:30  */
  assign i_control_fsm_n179 = i_control_fsm_adrx_mux_o; // (signal)
  /* mc8051_control_struc.vhd:148:30  */
  assign i_control_fsm_n180 = i_control_fsm_wrx_mux_o; // (signal)
  /* mc8051_control_struc.vhd:149:30  */
  assign i_control_fsm_n181 = i_control_fsm_data_mux_o; // (signal)
  /* mc8051_control_struc.vhd:150:30  */
  assign i_control_fsm_n182 = i_control_fsm_bdata_mux_o; // (signal)
  /* mc8051_control_struc.vhd:151:30  */
  assign i_control_fsm_n183 = i_control_fsm_regs_wr_en_o; // (signal)
  /* mc8051_control_struc.vhd:152:30  */
  assign i_control_fsm_n184 = i_control_fsm_help_en_o; // (signal)
  /* mc8051_control_struc.vhd:153:30  */
  assign i_control_fsm_n185 = i_control_fsm_help16_en_o; // (signal)
  /* mc8051_control_struc.vhd:154:30  */
  assign i_control_fsm_n186 = i_control_fsm_helpb_en_o; // (signal)
  /* mc8051_control_struc.vhd:155:30  */
  assign i_control_fsm_n187 = i_control_fsm_inthigh_en_o; // (signal)
  /* mc8051_control_struc.vhd:156:30  */
  assign i_control_fsm_n188 = i_control_fsm_intlow_en_o; // (signal)
  /* mc8051_control_struc.vhd:157:30  */
  assign i_control_fsm_n189 = i_control_fsm_intpre2_en_o; // (signal)
  /* mc8051_control_struc.vhd:158:30  */
  assign i_control_fsm_n190 = i_control_fsm_inthigh_d_o; // (signal)
  /* mc8051_control_struc.vhd:159:30  */
  assign i_control_fsm_n191 = i_control_fsm_intlow_d_o; // (signal)
  /* mc8051_control_struc.vhd:160:30  */
  assign i_control_fsm_n192 = i_control_fsm_intpre2_d_o; // (signal)
  /* mc8051_control_struc.vhd:161:31  */
  assign i_control_fsm_n193 = i_control_fsm_ext0isr_d_o; // (signal)
  /* mc8051_control_struc.vhd:162:31  */
  assign i_control_fsm_n194 = i_control_fsm_ext1isr_d_o; // (signal)
  /* mc8051_control_struc.vhd:163:31  */
  assign i_control_fsm_n195 = i_control_fsm_ext0isrh_d_o; // (signal)
  /* mc8051_control_struc.vhd:164:31  */
  assign i_control_fsm_n196 = i_control_fsm_ext1isrh_d_o; // (signal)
  /* mc8051_control_struc.vhd:165:31  */
  assign i_control_fsm_n197 = i_control_fsm_ext0isr_en_o; // (signal)
  /* mc8051_control_struc.vhd:166:31  */
  assign i_control_fsm_n198 = i_control_fsm_ext1isr_en_o; // (signal)
  /* mc8051_control_struc.vhd:167:31  */
  assign i_control_fsm_n199 = i_control_fsm_ext0isrh_en_o; // (signal)
  /* mc8051_control_struc.vhd:168:31  */
  assign i_control_fsm_n200 = i_control_fsm_ext1isrh_en_o; // (signal)
  /* mc8051_control_struc.vhd:121:3  */
  control_fsm i_control_fsm (
    .state_i(state),
    .help_i(s_help),
    .bit_data_i(s_bit_data),
    .aludata_i(aludata_i),
    .command_i(s_command),
    .inthigh_i(s_inthigh),
    .intlow_i(s_intlow),
    .intpre_i(s_intpre),
    .intpre2_i(s_intpre2),
    .intblock_i(s_intblock),
    .ti_i(s_ti),
    .ri_i(s_ri),
    .ie0_i(s_ie0),
    .ie1_i(s_ie1),
    .tf0_i(s_tf0),
    .tf1_i(s_tf1),
    .acc(acc),
    .psw(psw),
    .ie(ie),
    .ip(ip),
    .alu_cmd_o(i_control_fsm_alu_cmd_o),
    .pc_inc_en_o(i_control_fsm_pc_inc_en_o),
    .nextstate_o(i_control_fsm_nextstate_o),
    .adr_mux_o(i_control_fsm_adr_mux_o),
    .adrx_mux_o(i_control_fsm_adrx_mux_o),
    .wrx_mux_o(i_control_fsm_wrx_mux_o),
    .data_mux_o(i_control_fsm_data_mux_o),
    .bdata_mux_o(i_control_fsm_bdata_mux_o),
    .regs_wr_en_o(i_control_fsm_regs_wr_en_o),
    .help_en_o(i_control_fsm_help_en_o),
    .help16_en_o(i_control_fsm_help16_en_o),
    .helpb_en_o(i_control_fsm_helpb_en_o),
    .inthigh_en_o(i_control_fsm_inthigh_en_o),
    .intlow_en_o(i_control_fsm_intlow_en_o),
    .intpre2_en_o(i_control_fsm_intpre2_en_o),
    .inthigh_d_o(i_control_fsm_inthigh_d_o),
    .intlow_d_o(i_control_fsm_intlow_d_o),
    .intpre2_d_o(i_control_fsm_intpre2_d_o),
    .ext0isr_d_o(i_control_fsm_ext0isr_d_o),
    .ext1isr_d_o(i_control_fsm_ext1isr_d_o),
    .ext0isrh_d_o(i_control_fsm_ext0isrh_d_o),
    .ext1isrh_d_o(i_control_fsm_ext1isrh_d_o),
    .ext0isr_en_o(i_control_fsm_ext0isr_en_o),
    .ext1isr_en_o(i_control_fsm_ext1isr_en_o),
    .ext0isrh_en_o(i_control_fsm_ext0isrh_en_o),
    .ext1isrh_en_o(i_control_fsm_ext1isrh_en_o));
  /* mc8051_control_struc.vhd:172:32  */
  assign i_control_mem_n253 = i_control_mem_pc_o; // (signal)
  /* mc8051_control_struc.vhd:174:32  */
  assign i_control_mem_n254 = i_control_mem_ram_data_o; // (signal)
  /* mc8051_control_struc.vhd:176:32  */
  assign i_control_mem_n255 = i_control_mem_ram_adr_o; // (signal)
  /* mc8051_control_struc.vhd:177:32  */
  assign i_control_mem_n256 = i_control_mem_reg_data_o; // (signal)
  /* mc8051_control_struc.vhd:178:32  */
  assign i_control_mem_n257 = i_control_mem_ram_wr_o; // (signal)
  /* mc8051_control_struc.vhd:179:32  */
  assign i_control_mem_n258 = i_control_mem_cy_o; // (signal)
  /* mc8051_control_struc.vhd:180:32  */
  assign i_control_mem_n259 = i_control_mem_ov_o; // (signal)
  /* mc8051_control_struc.vhd:181:32  */
  assign i_control_mem_n260 = i_control_mem_ram_en_o; // (signal)
  /* mc8051_control_struc.vhd:184:32  */
  assign i_control_mem_n261 = i_control_mem_acc_o; // (signal)
  /* mc8051_control_struc.vhd:196:32  */
  assign i_control_mem_n262 = i_control_mem_p0_o; // (signal)
  /* mc8051_control_struc.vhd:197:32  */
  assign i_control_mem_n263 = i_control_mem_p1_o; // (signal)
  /* mc8051_control_struc.vhd:198:32  */
  assign i_control_mem_n264 = i_control_mem_p2_o; // (signal)
  /* mc8051_control_struc.vhd:199:32  */
  assign i_control_mem_n265 = i_control_mem_p3_o; // (signal)
  /* mc8051_control_struc.vhd:200:32  */
  assign i_control_mem_n266 = i_control_mem_all_trans_o; // (signal)
  /* mc8051_control_struc.vhd:201:32  */
  assign i_control_mem_n267 = i_control_mem_all_scon_o; // (signal)
  /* mc8051_control_struc.vhd:202:32  */
  assign i_control_mem_n268 = i_control_mem_all_sbuf_o; // (signal)
  /* mc8051_control_struc.vhd:203:32  */
  assign i_control_mem_n269 = i_control_mem_all_smod_o; // (signal)
  /* mc8051_control_struc.vhd:206:32  */
  assign i_control_mem_n270 = i_control_mem_all_tcon_tr0_o; // (signal)
  /* mc8051_control_struc.vhd:207:32  */
  assign i_control_mem_n271 = i_control_mem_all_tcon_tr1_o; // (signal)
  /* mc8051_control_struc.vhd:208:32  */
  assign i_control_mem_n272 = i_control_mem_all_tmod_o; // (signal)
  /* mc8051_control_struc.vhd:209:32  */
  assign i_control_mem_n273 = i_control_mem_all_reload_o; // (signal)
  /* mc8051_control_struc.vhd:210:32  */
  assign i_control_mem_n274 = i_control_mem_all_wt_o; // (signal)
  /* mc8051_control_struc.vhd:211:32  */
  assign i_control_mem_n275 = i_control_mem_all_wt_en_o; // (signal)
  /* mc8051_control_struc.vhd:219:28  */
  assign i_control_mem_n276 = i_control_mem_state_o; // (signal)
  /* mc8051_control_struc.vhd:220:28  */
  assign i_control_mem_n277 = i_control_mem_help_o; // (signal)
  /* mc8051_control_struc.vhd:221:28  */
  assign i_control_mem_n278 = i_control_mem_bit_data_o; // (signal)
  /* mc8051_control_struc.vhd:222:28  */
  assign i_control_mem_n279 = i_control_mem_command_o; // (signal)
  /* mc8051_control_struc.vhd:223:28  */
  assign i_control_mem_n280 = i_control_mem_inthigh_o; // (signal)
  /* mc8051_control_struc.vhd:224:28  */
  assign i_control_mem_n281 = i_control_mem_intlow_o; // (signal)
  /* mc8051_control_struc.vhd:225:28  */
  assign i_control_mem_n282 = i_control_mem_intpre_o; // (signal)
  /* mc8051_control_struc.vhd:226:28  */
  assign i_control_mem_n283 = i_control_mem_intpre2_o; // (signal)
  /* mc8051_control_struc.vhd:227:28  */
  assign i_control_mem_n284 = i_control_mem_intblock_o; // (signal)
  /* mc8051_control_struc.vhd:228:28  */
  assign i_control_mem_n285 = i_control_mem_ti_o; // (signal)
  /* mc8051_control_struc.vhd:229:28  */
  assign i_control_mem_n286 = i_control_mem_ri_o; // (signal)
  /* mc8051_control_struc.vhd:230:28  */
  assign i_control_mem_n287 = i_control_mem_ie0_o; // (signal)
  /* mc8051_control_struc.vhd:231:28  */
  assign i_control_mem_n288 = i_control_mem_ie1_o; // (signal)
  /* mc8051_control_struc.vhd:232:28  */
  assign i_control_mem_n289 = i_control_mem_tf0_o; // (signal)
  /* mc8051_control_struc.vhd:233:28  */
  assign i_control_mem_n290 = i_control_mem_tf1_o; // (signal)
  /* mc8051_control_struc.vhd:234:28  */
  assign i_control_mem_n291 = i_control_mem_psw_o; // (signal)
  /* mc8051_control_struc.vhd:235:28  */
  assign i_control_mem_n292 = i_control_mem_ie_o; // (signal)
  /* mc8051_control_struc.vhd:236:28  */
  assign i_control_mem_n293 = i_control_mem_ip_o; // (signal)
  /* mc8051_control_struc.vhd:237:28  */
  assign i_control_mem_n294 = i_control_mem_adrx_o; // (signal)
  /* mc8051_control_struc.vhd:238:28  */
  assign i_control_mem_n295 = i_control_mem_datax_o; // (signal)
  /* mc8051_control_struc.vhd:240:28  */
  assign i_control_mem_n296 = i_control_mem_memx_o; // (signal)
  /* mc8051_control_struc.vhd:239:28  */
  assign i_control_mem_n297 = i_control_mem_wrx_o; // (signal)
  /* mc8051_control_struc.vhd:171:3  */
  control_mem i_control_mem (
    .rom_data_i(rom_data_i),
    .ram_data_i(ram_data_i),
    .aludata_i(aludata_i),
    .aludatb_i(aludatb_i),
    .new_cy_i(new_cy_i),
    .new_ov_i(new_ov_i),
    .reset(reset),
    .clk(clk),
    .cen(cen),
    .int0_i(int0_i),
    .int1_i(int1_i),
    .p0_i(p0_i),
    .p1_i(p1_i),
    .p2_i(p2_i),
    .p3_i(p3_i),
    .all_scon_i(all_scon_i),
    .all_sbuf_i(all_sbuf_i),
    .all_tf0_i(all_tf0_i),
    .all_tf1_i(all_tf1_i),
    .all_tl0_i(all_tl0_i),
    .all_tl1_i(all_tl1_i),
    .all_th0_i(all_th0_i),
    .all_th1_i(all_th1_i),
    .datax_i(datax_i),
    .pc_inc_en_i(s_pc_inc_en),
    .nextstate_i(s_nextstate),
    .adr_mux_i(s_adr_mux),
    .adrx_mux_i(s_adrx_mux),
    .wrx_mux_i(s_wrx_mux),
    .data_mux_i(s_data_mux),
    .bdata_mux_i(s_bdata_mux),
    .regs_wr_en_i(s_regs_wr_en),
    .help_en_i(s_help_en),
    .help16_en_i(s_help16_en),
    .helpb_en_i(s_helpb_en),
    .inthigh_en_i(s_inthigh_en),
    .intlow_en_i(s_intlow_en),
    .intpre2_en_i(s_intpre2_en),
    .inthigh_d_i(s_inthigh_d),
    .intlow_d_i(s_intlow_d),
    .intpre2_d_i(s_intpre2_d),
    .ext0isr_d_i(s_ext0isr_d),
    .ext1isr_d_i(s_ext1isr_d),
    .ext0isrh_d_i(s_ext0isrh_d),
    .ext1isrh_d_i(s_ext1isrh_d),
    .ext0isr_en_i(s_ext0isr_en),
    .ext1isr_en_i(s_ext1isr_en),
    .ext0isrh_en_i(s_ext0isrh_en),
    .ext1isrh_en_i(s_ext1isrh_en),
    .pc_o(i_control_mem_pc_o),
    .ram_data_o(i_control_mem_ram_data_o),
    .ram_adr_o(i_control_mem_ram_adr_o),
    .reg_data_o(i_control_mem_reg_data_o),
    .ram_wr_o(i_control_mem_ram_wr_o),
    .cy_o(i_control_mem_cy_o),
    .ov_o(i_control_mem_ov_o),
    .ram_en_o(i_control_mem_ram_en_o),
    .acc_o(i_control_mem_acc_o),
    .p0_o(i_control_mem_p0_o),
    .p1_o(i_control_mem_p1_o),
    .p2_o(i_control_mem_p2_o),
    .p3_o(i_control_mem_p3_o),
    .all_trans_o(i_control_mem_all_trans_o),
    .all_scon_o(i_control_mem_all_scon_o),
    .all_sbuf_o(i_control_mem_all_sbuf_o),
    .all_smod_o(i_control_mem_all_smod_o),
    .all_tcon_tr0_o(i_control_mem_all_tcon_tr0_o),
    .all_tcon_tr1_o(i_control_mem_all_tcon_tr1_o),
    .all_tmod_o(i_control_mem_all_tmod_o),
    .all_reload_o(i_control_mem_all_reload_o),
    .all_wt_o(i_control_mem_all_wt_o),
    .all_wt_en_o(i_control_mem_all_wt_en_o),
    .state_o(i_control_mem_state_o),
    .help_o(i_control_mem_help_o),
    .bit_data_o(i_control_mem_bit_data_o),
    .command_o(i_control_mem_command_o),
    .inthigh_o(i_control_mem_inthigh_o),
    .intlow_o(i_control_mem_intlow_o),
    .intpre_o(i_control_mem_intpre_o),
    .intpre2_o(i_control_mem_intpre2_o),
    .intblock_o(i_control_mem_intblock_o),
    .ti_o(i_control_mem_ti_o),
    .ri_o(i_control_mem_ri_o),
    .ie0_o(i_control_mem_ie0_o),
    .ie1_o(i_control_mem_ie1_o),
    .tf0_o(i_control_mem_tf0_o),
    .tf1_o(i_control_mem_tf1_o),
    .psw_o(i_control_mem_psw_o),
    .ie_o(i_control_mem_ie_o),
    .ip_o(i_control_mem_ip_o),
    .adrx_o(i_control_mem_adrx_o),
    .datax_o(i_control_mem_datax_o),
    .wrx_o(i_control_mem_wrx_o),
    .memx_o(i_control_mem_memx_o));
endmodule

module mc8051_core
  (input  clk,
   input  cen,
   input  reset,
   input  [7:0] rom_data_i,
   input  [7:0] ram_data_i,
   input  int0_i,
   input  int1_i,
   input  all_t0_i,
   input  all_t1_i,
   input  all_rxd_i,
   input  [7:0] p0_i,
   input  [7:0] p1_i,
   input  [7:0] p2_i,
   input  [7:0] p3_i,
   input  [7:0] datax_i,
   output [7:0] p0_o,
   output [7:0] p1_o,
   output [7:0] p2_o,
   output [7:0] p3_o,
   output all_rxd_o,
   output all_txd_o,
   output all_rxdwr_o,
   output [15:0] rom_adr_o,
   output [7:0] ram_data_o,
   output [6:0] ram_adr_o,
   output ram_wr_o,
   output ram_en_o,
   output [7:0] datax_o,
   output [15:0] adrx_o,
   output memx_o,
   output wrx_o);
  wire [7:0] s_reg_data;
  wire [1:0] s_cy;
  wire s_ov;
  wire [5:0] s_alu_cmd;
  wire [7:0] s_alu_data0;
  wire [7:0] s_alu_data1;
  wire [7:0] s_acc;
  wire [1:0] s_cyb;
  wire s_ovb;
  wire s_all_trans;
  wire [5:0] s_all_scon;
  wire [7:0] s_all_sbuf;
  wire s_all_smod;
  wire [2:0] s_all_scon_out;
  wire [7:0] s_all_sbuf_out;
  wire s_all_tcon_tr0;
  wire s_all_tcon_tr1;
  wire [7:0] s_all_tmod;
  wire [7:0] s_all_reload;
  wire [1:0] s_all_wt;
  wire s_all_wt_en;
  wire s_all_tf0;
  wire s_all_tf1;
  wire [7:0] s_all_tl0;
  wire [7:0] s_all_th0;
  wire [7:0] s_all_tl1;
  wire [7:0] s_all_th1;
  wire [15:0] i_mc8051_control_n16;
  wire [7:0] i_mc8051_control_n17;
  wire [6:0] i_mc8051_control_n18;
  wire [7:0] i_mc8051_control_n19;
  wire i_mc8051_control_n20;
  wire [1:0] i_mc8051_control_n21;
  wire i_mc8051_control_n22;
  wire i_mc8051_control_n23;
  wire [5:0] i_mc8051_control_n24;
  wire [7:0] i_mc8051_control_n25;
  wire [7:0] i_mc8051_control_n26;
  wire [15:0] i_mc8051_control_n27;
  wire i_mc8051_control_n28;
  wire i_mc8051_control_n29;
  wire [7:0] i_mc8051_control_n30;
  wire [7:0] i_mc8051_control_n31;
  wire [7:0] i_mc8051_control_n32;
  wire [7:0] i_mc8051_control_n33;
  wire i_mc8051_control_n34;
  wire [5:0] i_mc8051_control_n35;
  wire [7:0] i_mc8051_control_n36;
  wire i_mc8051_control_n37;
  wire i_mc8051_control_n38;
  wire i_mc8051_control_n39;
  wire [7:0] i_mc8051_control_n40;
  wire [7:0] i_mc8051_control_n41;
  wire [1:0] i_mc8051_control_n42;
  wire i_mc8051_control_n43;
  wire [15:0] i_mc8051_control_pc_o;
  wire [7:0] i_mc8051_control_ram_data_o;
  wire [6:0] i_mc8051_control_ram_adr_o;
  wire [7:0] i_mc8051_control_reg_data_o;
  wire i_mc8051_control_ram_wr_o;
  wire [1:0] i_mc8051_control_cy_o;
  wire i_mc8051_control_ov_o;
  wire i_mc8051_control_ram_en_o;
  wire [5:0] i_mc8051_control_alu_cmd_o;
  wire [7:0] i_mc8051_control_acc_o;
  wire [7:0] i_mc8051_control_datax_o;
  wire [15:0] i_mc8051_control_adrx_o;
  wire i_mc8051_control_wrx_o;
  wire i_mc8051_control_memx_o;
  wire [7:0] i_mc8051_control_p0_o;
  wire [7:0] i_mc8051_control_p1_o;
  wire [7:0] i_mc8051_control_p2_o;
  wire [7:0] i_mc8051_control_p3_o;
  wire i_mc8051_control_all_trans_o;
  wire [5:0] i_mc8051_control_all_scon_o;
  wire [7:0] i_mc8051_control_all_sbuf_o;
  wire i_mc8051_control_all_smod_o;
  wire i_mc8051_control_all_tcon_tr0_o;
  wire i_mc8051_control_all_tcon_tr1_o;
  wire [7:0] i_mc8051_control_all_tmod_o;
  wire [7:0] i_mc8051_control_all_reload_o;
  wire [1:0] i_mc8051_control_all_wt_o;
  wire i_mc8051_control_all_wt_en_o;
  wire [1:0] i_mc8051_alu_n100;
  wire i_mc8051_alu_n101;
  wire [7:0] i_mc8051_alu_n102;
  wire [7:0] i_mc8051_alu_n103;
  wire [1:0] i_mc8051_alu_new_cy_o;
  wire i_mc8051_alu_new_ov_o;
  wire [7:0] i_mc8051_alu_result_a_o;
  wire [7:0] i_mc8051_alu_result_b_o;
  wire [7:0] gen_mc8051_siu_n1_i_mc8051_siu_n112;
  wire [2:0] gen_mc8051_siu_n1_i_mc8051_siu_n113;
  wire gen_mc8051_siu_n1_i_mc8051_siu_n114;
  wire gen_mc8051_siu_n1_i_mc8051_siu_n115;
  wire gen_mc8051_siu_n1_i_mc8051_siu_n116;
  wire [7:0] gen_mc8051_siu_n1_i_mc8051_siu_sbuf_o;
  wire [2:0] gen_mc8051_siu_n1_i_mc8051_siu_scon_o;
  wire gen_mc8051_siu_n1_i_mc8051_siu_rxdwr_o;
  wire gen_mc8051_siu_n1_i_mc8051_siu_rxd_o;
  wire gen_mc8051_siu_n1_i_mc8051_siu_txd_o;
  wire [7:0] gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n127;
  wire [7:0] gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n128;
  wire [7:0] gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n129;
  wire [7:0] gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n130;
  wire gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n131;
  wire gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n132;
  wire [7:0] gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_th0_o;
  wire [7:0] gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tl0_o;
  wire [7:0] gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_th1_o;
  wire [7:0] gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tl1_o;
  wire gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tf0_o;
  wire gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tf1_o;
  assign p0_o = i_mc8051_control_n30;
  assign p1_o = i_mc8051_control_n31;
  assign p2_o = i_mc8051_control_n32;
  assign p3_o = i_mc8051_control_n33;
  assign all_rxd_o = gen_mc8051_siu_n1_i_mc8051_siu_n115;
  assign all_txd_o = gen_mc8051_siu_n1_i_mc8051_siu_n116;
  assign all_rxdwr_o = gen_mc8051_siu_n1_i_mc8051_siu_n114;
  assign rom_adr_o = i_mc8051_control_n16;
  assign ram_data_o = i_mc8051_control_n17;
  assign ram_adr_o = i_mc8051_control_n18;
  assign ram_wr_o = i_mc8051_control_n20;
  assign ram_en_o = i_mc8051_control_n23;
  assign datax_o = i_mc8051_control_n26;
  assign adrx_o = i_mc8051_control_n27;
  assign memx_o = i_mc8051_control_n28;
  assign wrx_o = i_mc8051_control_n29;
  /* mc8051_core_struc.vhd:71:10  */
  assign s_reg_data = i_mc8051_control_n19; // (signal)
  /* mc8051_core_struc.vhd:72:10  */
  assign s_cy = i_mc8051_control_n21; // (signal)
  /* mc8051_core_struc.vhd:73:10  */
  assign s_ov = i_mc8051_control_n22; // (signal)
  /* mc8051_core_struc.vhd:74:10  */
  assign s_alu_cmd = i_mc8051_control_n24; // (signal)
  /* mc8051_core_struc.vhd:75:10  */
  assign s_alu_data0 = i_mc8051_alu_n102; // (signal)
  /* mc8051_core_struc.vhd:76:10  */
  assign s_alu_data1 = i_mc8051_alu_n103; // (signal)
  /* mc8051_core_struc.vhd:77:10  */
  assign s_acc = i_mc8051_control_n25; // (signal)
  /* mc8051_core_struc.vhd:78:10  */
  assign s_cyb = i_mc8051_alu_n100; // (signal)
  /* mc8051_core_struc.vhd:79:10  */
  assign s_ovb = i_mc8051_alu_n101; // (signal)
  /* mc8051_core_struc.vhd:185:41  */
  assign s_all_trans = i_mc8051_control_n34; // (signal)
  /* mc8051_core_struc.vhd:187:40  */
  assign s_all_scon = i_mc8051_control_n35; // (signal)
  /* mc8051_core_struc.vhd:188:40  */
  assign s_all_sbuf = i_mc8051_control_n36; // (signal)
  /* mc8051_core_struc.vhd:189:40  */
  assign s_all_smod = i_mc8051_control_n37; // (signal)
  /* mc8051_core_struc.vhd:89:10  */
  assign s_all_scon_out = gen_mc8051_siu_n1_i_mc8051_siu_n113; // (signal)
  /* mc8051_core_struc.vhd:90:10  */
  assign s_all_sbuf_out = gen_mc8051_siu_n1_i_mc8051_siu_n112; // (signal)
  /* mc8051_core_struc.vhd:209:45  */
  assign s_all_tcon_tr0 = i_mc8051_control_n38; // (signal)
  /* mc8051_core_struc.vhd:210:45  */
  assign s_all_tcon_tr1 = i_mc8051_control_n39; // (signal)
  /* mc8051_core_struc.vhd:208:41  */
  assign s_all_tmod = i_mc8051_control_n40; // (signal)
  /* mc8051_core_struc.vhd:211:43  */
  assign s_all_reload = i_mc8051_control_n41; // (signal)
  /* mc8051_core_struc.vhd:213:39  */
  assign s_all_wt = i_mc8051_control_n42; // (signal)
  /* mc8051_core_struc.vhd:212:42  */
  assign s_all_wt_en = i_mc8051_control_n43; // (signal)
  /* mc8051_core_struc.vhd:100:10  */
  assign s_all_tf0 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n131; // (signal)
  /* mc8051_core_struc.vhd:184:39  */
  assign s_all_tf1 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n132; // (signal)
  /* mc8051_core_struc.vhd:102:10  */
  assign s_all_tl0 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n128; // (signal)
  /* mc8051_core_struc.vhd:103:10  */
  assign s_all_th0 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n127; // (signal)
  /* mc8051_core_struc.vhd:104:10  */
  assign s_all_tl1 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n130; // (signal)
  /* mc8051_core_struc.vhd:105:10  */
  assign s_all_th1 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n129; // (signal)
  /* mc8051_core_struc.vhd:110:32  */
  assign i_mc8051_control_n16 = i_mc8051_control_pc_o; // (signal)
  /* mc8051_core_struc.vhd:112:32  */
  assign i_mc8051_control_n17 = i_mc8051_control_ram_data_o; // (signal)
  /* mc8051_core_struc.vhd:114:32  */
  assign i_mc8051_control_n18 = i_mc8051_control_ram_adr_o; // (signal)
  /* mc8051_core_struc.vhd:115:32  */
  assign i_mc8051_control_n19 = i_mc8051_control_reg_data_o; // (signal)
  /* mc8051_core_struc.vhd:116:32  */
  assign i_mc8051_control_n20 = i_mc8051_control_ram_wr_o; // (signal)
  /* mc8051_core_struc.vhd:117:32  */
  assign i_mc8051_control_n21 = i_mc8051_control_cy_o; // (signal)
  /* mc8051_core_struc.vhd:118:32  */
  assign i_mc8051_control_n22 = i_mc8051_control_ov_o; // (signal)
  /* mc8051_core_struc.vhd:119:32  */
  assign i_mc8051_control_n23 = i_mc8051_control_ram_en_o; // (signal)
  /* mc8051_core_struc.vhd:120:32  */
  assign i_mc8051_control_n24 = i_mc8051_control_alu_cmd_o; // (signal)
  /* mc8051_core_struc.vhd:123:32  */
  assign i_mc8051_control_n25 = i_mc8051_control_acc_o; // (signal)
  /* mc8051_core_struc.vhd:158:32  */
  assign i_mc8051_control_n26 = i_mc8051_control_datax_o; // (signal)
  /* mc8051_core_struc.vhd:157:32  */
  assign i_mc8051_control_n27 = i_mc8051_control_adrx_o; // (signal)
  /* mc8051_core_struc.vhd:160:32  */
  assign i_mc8051_control_n28 = i_mc8051_control_memx_o; // (signal)
  /* mc8051_core_struc.vhd:159:32  */
  assign i_mc8051_control_n29 = i_mc8051_control_wrx_o; // (signal)
  /* mc8051_core_struc.vhd:135:32  */
  assign i_mc8051_control_n30 = i_mc8051_control_p0_o; // (signal)
  /* mc8051_core_struc.vhd:136:32  */
  assign i_mc8051_control_n31 = i_mc8051_control_p1_o; // (signal)
  /* mc8051_core_struc.vhd:137:32  */
  assign i_mc8051_control_n32 = i_mc8051_control_p2_o; // (signal)
  /* mc8051_core_struc.vhd:138:32  */
  assign i_mc8051_control_n33 = i_mc8051_control_p3_o; // (signal)
  /* mc8051_core_struc.vhd:139:32  */
  assign i_mc8051_control_n34 = i_mc8051_control_all_trans_o; // (signal)
  /* mc8051_core_struc.vhd:140:32  */
  assign i_mc8051_control_n35 = i_mc8051_control_all_scon_o; // (signal)
  /* mc8051_core_struc.vhd:141:32  */
  assign i_mc8051_control_n36 = i_mc8051_control_all_sbuf_o; // (signal)
  /* mc8051_core_struc.vhd:142:32  */
  assign i_mc8051_control_n37 = i_mc8051_control_all_smod_o; // (signal)
  /* mc8051_core_struc.vhd:145:32  */
  assign i_mc8051_control_n38 = i_mc8051_control_all_tcon_tr0_o; // (signal)
  /* mc8051_core_struc.vhd:146:32  */
  assign i_mc8051_control_n39 = i_mc8051_control_all_tcon_tr1_o; // (signal)
  /* mc8051_core_struc.vhd:147:32  */
  assign i_mc8051_control_n40 = i_mc8051_control_all_tmod_o; // (signal)
  /* mc8051_core_struc.vhd:148:32  */
  assign i_mc8051_control_n41 = i_mc8051_control_all_reload_o; // (signal)
  /* mc8051_core_struc.vhd:149:32  */
  assign i_mc8051_control_n42 = i_mc8051_control_all_wt_o; // (signal)
  /* mc8051_core_struc.vhd:150:32  */
  assign i_mc8051_control_n43 = i_mc8051_control_all_wt_en_o; // (signal)
  /* mc8051_core_struc.vhd:109:3  */
  mc8051_control i_mc8051_control (
    .rom_data_i(rom_data_i),
    .ram_data_i(ram_data_i),
    .aludata_i(s_alu_data0),
    .aludatb_i(s_alu_data1),
    .new_cy_i(s_cyb),
    .new_ov_i(s_ovb),
    .reset(reset),
    .clk(clk),
    .cen(cen),
    .int0_i(int0_i),
    .int1_i(int1_i),
    .datax_i(datax_i),
    .p0_i(p0_i),
    .p1_i(p1_i),
    .p2_i(p2_i),
    .p3_i(p3_i),
    .all_scon_i(s_all_scon_out),
    .all_sbuf_i(s_all_sbuf_out),
    .all_tf0_i(s_all_tf0),
    .all_tf1_i(s_all_tf1),
    .all_tl0_i(s_all_tl0),
    .all_tl1_i(s_all_tl1),
    .all_th0_i(s_all_th0),
    .all_th1_i(s_all_th1),
    .pc_o(i_mc8051_control_pc_o),
    .ram_data_o(i_mc8051_control_ram_data_o),
    .ram_adr_o(i_mc8051_control_ram_adr_o),
    .reg_data_o(i_mc8051_control_reg_data_o),
    .ram_wr_o(i_mc8051_control_ram_wr_o),
    .cy_o(i_mc8051_control_cy_o),
    .ov_o(i_mc8051_control_ov_o),
    .ram_en_o(i_mc8051_control_ram_en_o),
    .alu_cmd_o(i_mc8051_control_alu_cmd_o),
    .acc_o(i_mc8051_control_acc_o),
    .datax_o(i_mc8051_control_datax_o),
    .adrx_o(i_mc8051_control_adrx_o),
    .wrx_o(i_mc8051_control_wrx_o),
    .memx_o(i_mc8051_control_memx_o),
    .p0_o(i_mc8051_control_p0_o),
    .p1_o(i_mc8051_control_p1_o),
    .p2_o(i_mc8051_control_p2_o),
    .p3_o(i_mc8051_control_p3_o),
    .all_trans_o(i_mc8051_control_all_trans_o),
    .all_scon_o(i_mc8051_control_all_scon_o),
    .all_sbuf_o(i_mc8051_control_all_sbuf_o),
    .all_smod_o(i_mc8051_control_all_smod_o),
    .all_tcon_tr0_o(i_mc8051_control_all_tcon_tr0_o),
    .all_tcon_tr1_o(i_mc8051_control_all_tcon_tr1_o),
    .all_tmod_o(i_mc8051_control_all_tmod_o),
    .all_reload_o(i_mc8051_control_all_reload_o),
    .all_wt_o(i_mc8051_control_all_wt_o),
    .all_wt_en_o(i_mc8051_control_all_wt_en_o));
  /* mc8051_core_struc.vhd:175:28  */
  assign i_mc8051_alu_n100 = i_mc8051_alu_new_cy_o; // (signal)
  /* mc8051_core_struc.vhd:176:28  */
  assign i_mc8051_alu_n101 = i_mc8051_alu_new_ov_o; // (signal)
  /* mc8051_core_struc.vhd:173:28  */
  assign i_mc8051_alu_n102 = i_mc8051_alu_result_a_o; // (signal)
  /* mc8051_core_struc.vhd:174:28  */
  assign i_mc8051_alu_n103 = i_mc8051_alu_result_b_o; // (signal)
  /* mc8051_core_struc.vhd:164:3  */
  mc8051_alu_8 i_mc8051_alu (
    .rom_data_i(rom_data_i),
    .ram_data_i(s_reg_data),
    .acc_i(s_acc),
    .cmd_i(s_alu_cmd),
    .cy_i(s_cy),
    .ov_i(s_ov),
    .new_cy_o(i_mc8051_alu_new_cy_o),
    .new_ov_o(i_mc8051_alu_new_ov_o),
    .result_a_o(i_mc8051_alu_result_a_o),
    .result_b_o(i_mc8051_alu_result_b_o));
  /* mc8051_core_struc.vhd:191:30  */
  assign gen_mc8051_siu_n1_i_mc8051_siu_n112 = gen_mc8051_siu_n1_i_mc8051_siu_sbuf_o; // (signal)
  /* mc8051_core_struc.vhd:192:30  */
  assign gen_mc8051_siu_n1_i_mc8051_siu_n113 = gen_mc8051_siu_n1_i_mc8051_siu_scon_o; // (signal)
  /* mc8051_core_struc.vhd:193:30  */
  assign gen_mc8051_siu_n1_i_mc8051_siu_n114 = gen_mc8051_siu_n1_i_mc8051_siu_rxdwr_o; // (signal)
  /* mc8051_core_struc.vhd:194:30  */
  assign gen_mc8051_siu_n1_i_mc8051_siu_n115 = gen_mc8051_siu_n1_i_mc8051_siu_rxd_o; // (signal)
  /* mc8051_core_struc.vhd:195:30  */
  assign gen_mc8051_siu_n1_i_mc8051_siu_n116 = gen_mc8051_siu_n1_i_mc8051_siu_txd_o; // (signal)
  /* mc8051_core_struc.vhd:180:5  */
  mc8051_siu gen_mc8051_siu_n1_i_mc8051_siu (
    .clk(clk),
    .cen(cen),
    .reset(reset),
    .tf_i(s_all_tf1),
    .trans_i(s_all_trans),
    .rxd_i(all_rxd_i),
    .scon_i(s_all_scon),
    .sbuf_i(s_all_sbuf),
    .smod_i(s_all_smod),
    .sbuf_o(gen_mc8051_siu_n1_i_mc8051_siu_sbuf_o),
    .scon_o(gen_mc8051_siu_n1_i_mc8051_siu_scon_o),
    .rxdwr_o(gen_mc8051_siu_n1_i_mc8051_siu_rxdwr_o),
    .rxd_o(gen_mc8051_siu_n1_i_mc8051_siu_rxd_o),
    .txd_o(gen_mc8051_siu_n1_i_mc8051_siu_txd_o));
  /* mc8051_core_struc.vhd:215:31  */
  assign gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n127 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_th0_o; // (signal)
  /* mc8051_core_struc.vhd:216:31  */
  assign gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n128 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tl0_o; // (signal)
  /* mc8051_core_struc.vhd:217:31  */
  assign gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n129 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_th1_o; // (signal)
  /* mc8051_core_struc.vhd:218:31  */
  assign gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n130 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tl1_o; // (signal)
  /* mc8051_core_struc.vhd:219:31  */
  assign gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n131 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tf0_o; // (signal)
  /* mc8051_core_struc.vhd:220:31  */
  assign gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_n132 = gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tf1_o; // (signal)
  /* mc8051_core_struc.vhd:200:5  */
  mc8051_tmrctr gen_mc8051_tmrctr_n1_i_mc8051_tmrctr (
    .clk(clk),
    .cen(cen),
    .reset(reset),
    .int0_i(int0_i),
    .int1_i(int1_i),
    .t0_i(all_t0_i),
    .t1_i(all_t1_i),
    .tmod_i(s_all_tmod),
    .tcon_tr0_i(s_all_tcon_tr0),
    .tcon_tr1_i(s_all_tcon_tr1),
    .reload_i(s_all_reload),
    .wt_en_i(s_all_wt_en),
    .wt_i(s_all_wt),
    .th0_o(gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_th0_o),
    .tl0_o(gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tl0_o),
    .th1_o(gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_th1_o),
    .tl1_o(gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tl1_o),
    .tf0_o(gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tf0_o),
    .tf1_o(gen_mc8051_tmrctr_n1_i_mc8051_tmrctr_tf1_o));
endmodule

